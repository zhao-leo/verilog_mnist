// MNIST手写数字识别模型 - Int8量化版本（串行计算架构）
// MNIST手写数字识别模型 - Int8量化版本（高度优化串行架构）
// 极致优化：3个隐藏神经元，24位累加器，最小化逻辑资源
// 网络结构: 784 → 3 → 10
// 输入: 28x28二值图像 (784位)
// 输出: 预测数字 (0-9)
// 时钟周期: ~2395 cycles
// ROM大小: 2395 bytes
// 优化目标: LUT < 6,272

module mnist_model(
    input wire clk,
    input wire rst,
    input wire [783:0] image_in,
    input wire start,
    output reg [3:0] digit_out,
    output reg valid
);

    // 紧凑状态机 (2位足够5个状态)
    localparam IDLE = 2'd0;
    localparam LAYER1 = 2'd1;
    localparam LAYER2 = 2'd2;
    localparam ARGMAX = 2'd3;

    reg [1:0] state;
    reg [3:0] neuron_idx;    // 神经元索引 (0-9)
    reg [9:0] input_idx;     // 输入索引 (0-783)
    reg layer1_done;         // Layer1计算完成标志

    // 24位累加器（减少寄存器使用）
    reg signed [23:0] accumulator;

    // 层输出存储（24位）
    reg signed [23:0] layer1_out [0:2];
    reg signed [23:0] layer2_out [0:9];

    // Argmax变量
    reg [3:0] max_idx;
    reg signed [23:0] max_val;

    // ROM: 权重和偏置 (2395字节)
    // 强制使用BRAM以节省LUT
    (* ram_style = "block" *)
    (* ramstyle = "M9K" *)
    (* syn_ramstyle = "block_ram" *)
    reg signed [7:0] weight_rom [0:2394];

    // 初始化ROM
    initial begin
        weight_rom[0] = 0;
        weight_rom[1] = -2;
        weight_rom[2] = -2;
        weight_rom[3] = 0;
        weight_rom[4] = 1;
        weight_rom[5] = 1;
        weight_rom[6] = 2;
        weight_rom[7] = 2;
        weight_rom[8] = 0;
        weight_rom[9] = 0;
        weight_rom[10] = 0;
        weight_rom[11] = 2;
        weight_rom[12] = 2;
        weight_rom[13] = -6;
        weight_rom[14] = -18;
        weight_rom[15] = 2;
        weight_rom[16] = 1;
        weight_rom[17] = -1;
        weight_rom[18] = 0;
        weight_rom[19] = -1;
        weight_rom[20] = 1;
        weight_rom[21] = 2;
        weight_rom[22] = -2;
        weight_rom[23] = 0;
        weight_rom[24] = -1;
        weight_rom[25] = 1;
        weight_rom[26] = -2;
        weight_rom[27] = -2;
        weight_rom[28] = -1;
        weight_rom[29] = 0;
        weight_rom[30] = 0;
        weight_rom[31] = -1;
        weight_rom[32] = -2;
        weight_rom[33] = -1;
        weight_rom[34] = 15;
        weight_rom[35] = 25;
        weight_rom[36] = 33;
        weight_rom[37] = 25;
        weight_rom[38] = 30;
        weight_rom[39] = 25;
        weight_rom[40] = 34;
        weight_rom[41] = 43;
        weight_rom[42] = -7;
        weight_rom[43] = 4;
        weight_rom[44] = -13;
        weight_rom[45] = 11;
        weight_rom[46] = 52;
        weight_rom[47] = 31;
        weight_rom[48] = 34;
        weight_rom[49] = 19;
        weight_rom[50] = 23;
        weight_rom[51] = 15;
        weight_rom[52] = -2;
        weight_rom[53] = -2;
        weight_rom[54] = 2;
        weight_rom[55] = -2;
        weight_rom[56] = 1;
        weight_rom[57] = 0;
        weight_rom[58] = 2;
        weight_rom[59] = 0;
        weight_rom[60] = 19;
        weight_rom[61] = -1;
        weight_rom[62] = 31;
        weight_rom[63] = 36;
        weight_rom[64] = 35;
        weight_rom[65] = 22;
        weight_rom[66] = 59;
        weight_rom[67] = 38;
        weight_rom[68] = 52;
        weight_rom[69] = 35;
        weight_rom[70] = 49;
        weight_rom[71] = 38;
        weight_rom[72] = 55;
        weight_rom[73] = 44;
        weight_rom[74] = 57;
        weight_rom[75] = 60;
        weight_rom[76] = 72;
        weight_rom[77] = 46;
        weight_rom[78] = 46;
        weight_rom[79] = 21;
        weight_rom[80] = 0;
        weight_rom[81] = -15;
        weight_rom[82] = -1;
        weight_rom[83] = 0;
        weight_rom[84] = 2;
        weight_rom[85] = 1;
        weight_rom[86] = 16;
        weight_rom[87] = -2;
        weight_rom[88] = -1;
        weight_rom[89] = -13;
        weight_rom[90] = 36;
        weight_rom[91] = 26;
        weight_rom[92] = 16;
        weight_rom[93] = 28;
        weight_rom[94] = 22;
        weight_rom[95] = 7;
        weight_rom[96] = 6;
        weight_rom[97] = 5;
        weight_rom[98] = 4;
        weight_rom[99] = 13;
        weight_rom[100] = 15;
        weight_rom[101] = 17;
        weight_rom[102] = 31;
        weight_rom[103] = 33;
        weight_rom[104] = 45;
        weight_rom[105] = 56;
        weight_rom[106] = 53;
        weight_rom[107] = 32;
        weight_rom[108] = 33;
        weight_rom[109] = -16;
        weight_rom[110] = 0;
        weight_rom[111] = -1;
        weight_rom[112] = 1;
        weight_rom[113] = 2;
        weight_rom[114] = -16;
        weight_rom[115] = 0;
        weight_rom[116] = 12;
        weight_rom[117] = 4;
        weight_rom[118] = 0;
        weight_rom[119] = 12;
        weight_rom[120] = 15;
        weight_rom[121] = 5;
        weight_rom[122] = 7;
        weight_rom[123] = 0;
        weight_rom[124] = -2;
        weight_rom[125] = 3;
        weight_rom[126] = 1;
        weight_rom[127] = -3;
        weight_rom[128] = -6;
        weight_rom[129] = -1;
        weight_rom[130] = -9;
        weight_rom[131] = -5;
        weight_rom[132] = -10;
        weight_rom[133] = -9;
        weight_rom[134] = -3;
        weight_rom[135] = 21;
        weight_rom[136] = 22;
        weight_rom[137] = -6;
        weight_rom[138] = -19;
        weight_rom[139] = 1;
        weight_rom[140] = 1;
        weight_rom[141] = -2;
        weight_rom[142] = 1;
        weight_rom[143] = -12;
        weight_rom[144] = -2;
        weight_rom[145] = -8;
        weight_rom[146] = 1;
        weight_rom[147] = 9;
        weight_rom[148] = 8;
        weight_rom[149] = 9;
        weight_rom[150] = 5;
        weight_rom[151] = -5;
        weight_rom[152] = 1;
        weight_rom[153] = -1;
        weight_rom[154] = 4;
        weight_rom[155] = -1;
        weight_rom[156] = 5;
        weight_rom[157] = 9;
        weight_rom[158] = 2;
        weight_rom[159] = 0;
        weight_rom[160] = -2;
        weight_rom[161] = -9;
        weight_rom[162] = -7;
        weight_rom[163] = -2;
        weight_rom[164] = 1;
        weight_rom[165] = 5;
        weight_rom[166] = -2;
        weight_rom[167] = -1;
        weight_rom[168] = 0;
        weight_rom[169] = 1;
        weight_rom[170] = -19;
        weight_rom[171] = -18;
        weight_rom[172] = 0;
        weight_rom[173] = 6;
        weight_rom[174] = -10;
        weight_rom[175] = 3;
        weight_rom[176] = 4;
        weight_rom[177] = 6;
        weight_rom[178] = 0;
        weight_rom[179] = -5;
        weight_rom[180] = -4;
        weight_rom[181] = -6;
        weight_rom[182] = -8;
        weight_rom[183] = -3;
        weight_rom[184] = -6;
        weight_rom[185] = 0;
        weight_rom[186] = -11;
        weight_rom[187] = -8;
        weight_rom[188] = -8;
        weight_rom[189] = -9;
        weight_rom[190] = -2;
        weight_rom[191] = 7;
        weight_rom[192] = 18;
        weight_rom[193] = 6;
        weight_rom[194] = -8;
        weight_rom[195] = 17;
        weight_rom[196] = 0;
        weight_rom[197] = -13;
        weight_rom[198] = -15;
        weight_rom[199] = -22;
        weight_rom[200] = -4;
        weight_rom[201] = -1;
        weight_rom[202] = -3;
        weight_rom[203] = 0;
        weight_rom[204] = 2;
        weight_rom[205] = -2;
        weight_rom[206] = 0;
        weight_rom[207] = -5;
        weight_rom[208] = -13;
        weight_rom[209] = -12;
        weight_rom[210] = -8;
        weight_rom[211] = -2;
        weight_rom[212] = -2;
        weight_rom[213] = -9;
        weight_rom[214] = -9;
        weight_rom[215] = -8;
        weight_rom[216] = -6;
        weight_rom[217] = -3;
        weight_rom[218] = 1;
        weight_rom[219] = 4;
        weight_rom[220] = 9;
        weight_rom[221] = 2;
        weight_rom[222] = -12;
        weight_rom[223] = -15;
        weight_rom[224] = 1;
        weight_rom[225] = -22;
        weight_rom[226] = -10;
        weight_rom[227] = -14;
        weight_rom[228] = -8;
        weight_rom[229] = -1;
        weight_rom[230] = -1;
        weight_rom[231] = -4;
        weight_rom[232] = -4;
        weight_rom[233] = 3;
        weight_rom[234] = -1;
        weight_rom[235] = -2;
        weight_rom[236] = -12;
        weight_rom[237] = -12;
        weight_rom[238] = -15;
        weight_rom[239] = -12;
        weight_rom[240] = -13;
        weight_rom[241] = -17;
        weight_rom[242] = -10;
        weight_rom[243] = -9;
        weight_rom[244] = -3;
        weight_rom[245] = 4;
        weight_rom[246] = 5;
        weight_rom[247] = -2;
        weight_rom[248] = 15;
        weight_rom[249] = 2;
        weight_rom[250] = -21;
        weight_rom[251] = 5;
        weight_rom[252] = -17;
        weight_rom[253] = -29;
        weight_rom[254] = -21;
        weight_rom[255] = -26;
        weight_rom[256] = -3;
        weight_rom[257] = -2;
        weight_rom[258] = 0;
        weight_rom[259] = -2;
        weight_rom[260] = -3;
        weight_rom[261] = 2;
        weight_rom[262] = 2;
        weight_rom[263] = -4;
        weight_rom[264] = -9;
        weight_rom[265] = -18;
        weight_rom[266] = -31;
        weight_rom[267] = -21;
        weight_rom[268] = -18;
        weight_rom[269] = -12;
        weight_rom[270] = -9;
        weight_rom[271] = -6;
        weight_rom[272] = 1;
        weight_rom[273] = 6;
        weight_rom[274] = 0;
        weight_rom[275] = 7;
        weight_rom[276] = 6;
        weight_rom[277] = 16;
        weight_rom[278] = -1;
        weight_rom[279] = -17;
        weight_rom[280] = -18;
        weight_rom[281] = -24;
        weight_rom[282] = -24;
        weight_rom[283] = -20;
        weight_rom[284] = 2;
        weight_rom[285] = -8;
        weight_rom[286] = 1;
        weight_rom[287] = 2;
        weight_rom[288] = 2;
        weight_rom[289] = 5;
        weight_rom[290] = 7;
        weight_rom[291] = 5;
        weight_rom[292] = 1;
        weight_rom[293] = -11;
        weight_rom[294] = -34;
        weight_rom[295] = -31;
        weight_rom[296] = -22;
        weight_rom[297] = -13;
        weight_rom[298] = -11;
        weight_rom[299] = -5;
        weight_rom[300] = -6;
        weight_rom[301] = -1;
        weight_rom[302] = -3;
        weight_rom[303] = -7;
        weight_rom[304] = -5;
        weight_rom[305] = 2;
        weight_rom[306] = 0;
        weight_rom[307] = -31;
        weight_rom[308] = -4;
        weight_rom[309] = -28;
        weight_rom[310] = -35;
        weight_rom[311] = -17;
        weight_rom[312] = -4;
        weight_rom[313] = 5;
        weight_rom[314] = 2;
        weight_rom[315] = -4;
        weight_rom[316] = 6;
        weight_rom[317] = 5;
        weight_rom[318] = 10;
        weight_rom[319] = 13;
        weight_rom[320] = 15;
        weight_rom[321] = -1;
        weight_rom[322] = -18;
        weight_rom[323] = -18;
        weight_rom[324] = 5;
        weight_rom[325] = 4;
        weight_rom[326] = -5;
        weight_rom[327] = 0;
        weight_rom[328] = -2;
        weight_rom[329] = 0;
        weight_rom[330] = -11;
        weight_rom[331] = -11;
        weight_rom[332] = -6;
        weight_rom[333] = -6;
        weight_rom[334] = -5;
        weight_rom[335] = 15;
        weight_rom[336] = -4;
        weight_rom[337] = -11;
        weight_rom[338] = -23;
        weight_rom[339] = -22;
        weight_rom[340] = 0;
        weight_rom[341] = -5;
        weight_rom[342] = 0;
        weight_rom[343] = 2;
        weight_rom[344] = 2;
        weight_rom[345] = 6;
        weight_rom[346] = 9;
        weight_rom[347] = 18;
        weight_rom[348] = 17;
        weight_rom[349] = 12;
        weight_rom[350] = -16;
        weight_rom[351] = 4;
        weight_rom[352] = 16;
        weight_rom[353] = 16;
        weight_rom[354] = 11;
        weight_rom[355] = 8;
        weight_rom[356] = 0;
        weight_rom[357] = -2;
        weight_rom[358] = -6;
        weight_rom[359] = 2;
        weight_rom[360] = 21;
        weight_rom[361] = -29;
        weight_rom[362] = -39;
        weight_rom[363] = 15;
        weight_rom[364] = 0;
        weight_rom[365] = 4;
        weight_rom[366] = -39;
        weight_rom[367] = -14;
        weight_rom[368] = -7;
        weight_rom[369] = 2;
        weight_rom[370] = 0;
        weight_rom[371] = 1;
        weight_rom[372] = 5;
        weight_rom[373] = 5;
        weight_rom[374] = 9;
        weight_rom[375] = 17;
        weight_rom[376] = 19;
        weight_rom[377] = 11;
        weight_rom[378] = 3;
        weight_rom[379] = 14;
        weight_rom[380] = 15;
        weight_rom[381] = 23;
        weight_rom[382] = 17;
        weight_rom[383] = 6;
        weight_rom[384] = 0;
        weight_rom[385] = 7;
        weight_rom[386] = -10;
        weight_rom[387] = 4;
        weight_rom[388] = 7;
        weight_rom[389] = -20;
        weight_rom[390] = -22;
        weight_rom[391] = -17;
        weight_rom[392] = -1;
        weight_rom[393] = -16;
        weight_rom[394] = -3;
        weight_rom[395] = 1;
        weight_rom[396] = 20;
        weight_rom[397] = 7;
        weight_rom[398] = 8;
        weight_rom[399] = 6;
        weight_rom[400] = 6;
        weight_rom[401] = 5;
        weight_rom[402] = 4;
        weight_rom[403] = 30;
        weight_rom[404] = 22;
        weight_rom[405] = 10;
        weight_rom[406] = 8;
        weight_rom[407] = 6;
        weight_rom[408] = 20;
        weight_rom[409] = 21;
        weight_rom[410] = 1;
        weight_rom[411] = -2;
        weight_rom[412] = -4;
        weight_rom[413] = -9;
        weight_rom[414] = -2;
        weight_rom[415] = -11;
        weight_rom[416] = 7;
        weight_rom[417] = -3;
        weight_rom[418] = -16;
        weight_rom[419] = 0;
        weight_rom[420] = -1;
        weight_rom[421] = -13;
        weight_rom[422] = -4;
        weight_rom[423] = 25;
        weight_rom[424] = -9;
        weight_rom[425] = 5;
        weight_rom[426] = 6;
        weight_rom[427] = 3;
        weight_rom[428] = 7;
        weight_rom[429] = 1;
        weight_rom[430] = 6;
        weight_rom[431] = 23;
        weight_rom[432] = 20;
        weight_rom[433] = 20;
        weight_rom[434] = 15;
        weight_rom[435] = 6;
        weight_rom[436] = 26;
        weight_rom[437] = 14;
        weight_rom[438] = -3;
        weight_rom[439] = -10;
        weight_rom[440] = -12;
        weight_rom[441] = -6;
        weight_rom[442] = -7;
        weight_rom[443] = -10;
        weight_rom[444] = -6;
        weight_rom[445] = 31;
        weight_rom[446] = 11;
        weight_rom[447] = 14;
        weight_rom[448] = 0;
        weight_rom[449] = -1;
        weight_rom[450] = -14;
        weight_rom[451] = 4;
        weight_rom[452] = -16;
        weight_rom[453] = 5;
        weight_rom[454] = 11;
        weight_rom[455] = 8;
        weight_rom[456] = 8;
        weight_rom[457] = 8;
        weight_rom[458] = 12;
        weight_rom[459] = 26;
        weight_rom[460] = 30;
        weight_rom[461] = 18;
        weight_rom[462] = 16;
        weight_rom[463] = 17;
        weight_rom[464] = 21;
        weight_rom[465] = 5;
        weight_rom[466] = -9;
        weight_rom[467] = -13;
        weight_rom[468] = -6;
        weight_rom[469] = -4;
        weight_rom[470] = -6;
        weight_rom[471] = -10;
        weight_rom[472] = 16;
        weight_rom[473] = 35;
        weight_rom[474] = -12;
        weight_rom[475] = -10;
        weight_rom[476] = 1;
        weight_rom[477] = -2;
        weight_rom[478] = 17;
        weight_rom[479] = -8;
        weight_rom[480] = -9;
        weight_rom[481] = -7;
        weight_rom[482] = -3;
        weight_rom[483] = 3;
        weight_rom[484] = 6;
        weight_rom[485] = 12;
        weight_rom[486] = 15;
        weight_rom[487] = 27;
        weight_rom[488] = 23;
        weight_rom[489] = 14;
        weight_rom[490] = 15;
        weight_rom[491] = 15;
        weight_rom[492] = 9;
        weight_rom[493] = -1;
        weight_rom[494] = -2;
        weight_rom[495] = -7;
        weight_rom[496] = -3;
        weight_rom[497] = -6;
        weight_rom[498] = -6;
        weight_rom[499] = -10;
        weight_rom[500] = 13;
        weight_rom[501] = 30;
        weight_rom[502] = 2;
        weight_rom[503] = 0;
        weight_rom[504] = -1;
        weight_rom[505] = 0;
        weight_rom[506] = -9;
        weight_rom[507] = 5;
        weight_rom[508] = -9;
        weight_rom[509] = 5;
        weight_rom[510] = -5;
        weight_rom[511] = 5;
        weight_rom[512] = 5;
        weight_rom[513] = 12;
        weight_rom[514] = 12;
        weight_rom[515] = 11;
        weight_rom[516] = 16;
        weight_rom[517] = 3;
        weight_rom[518] = 9;
        weight_rom[519] = 7;
        weight_rom[520] = 10;
        weight_rom[521] = 5;
        weight_rom[522] = 1;
        weight_rom[523] = 1;
        weight_rom[524] = 2;
        weight_rom[525] = -5;
        weight_rom[526] = -4;
        weight_rom[527] = 14;
        weight_rom[528] = 16;
        weight_rom[529] = 32;
        weight_rom[530] = 32;
        weight_rom[531] = -22;
        weight_rom[532] = 2;
        weight_rom[533] = -2;
        weight_rom[534] = -9;
        weight_rom[535] = -1;
        weight_rom[536] = -1;
        weight_rom[537] = -3;
        weight_rom[538] = 5;
        weight_rom[539] = 5;
        weight_rom[540] = 0;
        weight_rom[541] = 0;
        weight_rom[542] = 6;
        weight_rom[543] = 3;
        weight_rom[544] = -4;
        weight_rom[545] = 2;
        weight_rom[546] = 3;
        weight_rom[547] = 12;
        weight_rom[548] = 10;
        weight_rom[549] = 11;
        weight_rom[550] = 11;
        weight_rom[551] = 6;
        weight_rom[552] = 6;
        weight_rom[553] = 10;
        weight_rom[554] = 4;
        weight_rom[555] = 8;
        weight_rom[556] = 19;
        weight_rom[557] = 23;
        weight_rom[558] = 9;
        weight_rom[559] = -11;
        weight_rom[560] = 1;
        weight_rom[561] = -4;
        weight_rom[562] = 10;
        weight_rom[563] = 4;
        weight_rom[564] = 8;
        weight_rom[565] = 9;
        weight_rom[566] = -2;
        weight_rom[567] = 4;
        weight_rom[568] = 4;
        weight_rom[569] = 0;
        weight_rom[570] = -2;
        weight_rom[571] = -8;
        weight_rom[572] = -5;
        weight_rom[573] = -3;
        weight_rom[574] = -2;
        weight_rom[575] = 10;
        weight_rom[576] = 12;
        weight_rom[577] = 8;
        weight_rom[578] = 14;
        weight_rom[579] = 8;
        weight_rom[580] = 6;
        weight_rom[581] = 5;
        weight_rom[582] = 2;
        weight_rom[583] = 5;
        weight_rom[584] = 17;
        weight_rom[585] = 4;
        weight_rom[586] = 18;
        weight_rom[587] = 2;
        weight_rom[588] = 0;
        weight_rom[589] = 11;
        weight_rom[590] = 1;
        weight_rom[591] = 1;
        weight_rom[592] = 7;
        weight_rom[593] = 7;
        weight_rom[594] = 0;
        weight_rom[595] = 5;
        weight_rom[596] = -7;
        weight_rom[597] = -3;
        weight_rom[598] = -10;
        weight_rom[599] = -7;
        weight_rom[600] = -1;
        weight_rom[601] = -3;
        weight_rom[602] = 0;
        weight_rom[603] = -1;
        weight_rom[604] = 4;
        weight_rom[605] = 12;
        weight_rom[606] = 10;
        weight_rom[607] = 10;
        weight_rom[608] = 10;
        weight_rom[609] = 7;
        weight_rom[610] = 13;
        weight_rom[611] = 30;
        weight_rom[612] = 19;
        weight_rom[613] = -7;
        weight_rom[614] = 17;
        weight_rom[615] = 0;
        weight_rom[616] = 1;
        weight_rom[617] = 1;
        weight_rom[618] = -13;
        weight_rom[619] = 14;
        weight_rom[620] = 25;
        weight_rom[621] = 2;
        weight_rom[622] = -2;
        weight_rom[623] = -1;
        weight_rom[624] = -5;
        weight_rom[625] = -14;
        weight_rom[626] = -2;
        weight_rom[627] = -3;
        weight_rom[628] = 2;
        weight_rom[629] = 0;
        weight_rom[630] = -8;
        weight_rom[631] = -10;
        weight_rom[632] = -6;
        weight_rom[633] = -2;
        weight_rom[634] = 8;
        weight_rom[635] = 7;
        weight_rom[636] = 7;
        weight_rom[637] = 11;
        weight_rom[638] = 9;
        weight_rom[639] = 4;
        weight_rom[640] = 13;
        weight_rom[641] = -15;
        weight_rom[642] = -20;
        weight_rom[643] = 2;
        weight_rom[644] = -1;
        weight_rom[645] = 0;
        weight_rom[646] = -3;
        weight_rom[647] = 7;
        weight_rom[648] = -2;
        weight_rom[649] = -7;
        weight_rom[650] = -11;
        weight_rom[651] = -13;
        weight_rom[652] = 0;
        weight_rom[653] = -3;
        weight_rom[654] = -8;
        weight_rom[655] = 1;
        weight_rom[656] = -1;
        weight_rom[657] = 0;
        weight_rom[658] = -4;
        weight_rom[659] = -8;
        weight_rom[660] = -7;
        weight_rom[661] = -7;
        weight_rom[662] = 4;
        weight_rom[663] = 17;
        weight_rom[664] = 24;
        weight_rom[665] = 24;
        weight_rom[666] = 13;
        weight_rom[667] = 11;
        weight_rom[668] = -2;
        weight_rom[669] = 4;
        weight_rom[670] = -16;
        weight_rom[671] = -1;
        weight_rom[672] = 2;
        weight_rom[673] = -2;
        weight_rom[674] = 0;
        weight_rom[675] = -9;
        weight_rom[676] = -14;
        weight_rom[677] = -27;
        weight_rom[678] = -12;
        weight_rom[679] = -8;
        weight_rom[680] = 1;
        weight_rom[681] = 1;
        weight_rom[682] = 7;
        weight_rom[683] = 5;
        weight_rom[684] = 6;
        weight_rom[685] = 4;
        weight_rom[686] = 7;
        weight_rom[687] = 6;
        weight_rom[688] = 12;
        weight_rom[689] = 7;
        weight_rom[690] = 22;
        weight_rom[691] = 25;
        weight_rom[692] = 26;
        weight_rom[693] = 18;
        weight_rom[694] = 16;
        weight_rom[695] = 10;
        weight_rom[696] = -6;
        weight_rom[697] = 9;
        weight_rom[698] = -1;
        weight_rom[699] = 1;
        weight_rom[700] = -1;
        weight_rom[701] = 1;
        weight_rom[702] = -1;
        weight_rom[703] = 12;
        weight_rom[704] = -4;
        weight_rom[705] = -17;
        weight_rom[706] = -4;
        weight_rom[707] = 4;
        weight_rom[708] = -5;
        weight_rom[709] = -7;
        weight_rom[710] = 3;
        weight_rom[711] = -7;
        weight_rom[712] = -10;
        weight_rom[713] = -3;
        weight_rom[714] = 0;
        weight_rom[715] = -1;
        weight_rom[716] = 10;
        weight_rom[717] = 10;
        weight_rom[718] = 2;
        weight_rom[719] = -7;
        weight_rom[720] = 12;
        weight_rom[721] = -4;
        weight_rom[722] = 2;
        weight_rom[723] = -13;
        weight_rom[724] = -27;
        weight_rom[725] = 2;
        weight_rom[726] = 0;
        weight_rom[727] = -1;
        weight_rom[728] = 1;
        weight_rom[729] = -1;
        weight_rom[730] = 1;
        weight_rom[731] = -1;
        weight_rom[732] = 7;
        weight_rom[733] = -5;
        weight_rom[734] = 0;
        weight_rom[735] = -9;
        weight_rom[736] = -10;
        weight_rom[737] = -7;
        weight_rom[738] = -11;
        weight_rom[739] = -8;
        weight_rom[740] = 0;
        weight_rom[741] = -1;
        weight_rom[742] = -1;
        weight_rom[743] = 0;
        weight_rom[744] = -1;
        weight_rom[745] = -2;
        weight_rom[746] = 13;
        weight_rom[747] = 4;
        weight_rom[748] = 20;
        weight_rom[749] = 1;
        weight_rom[750] = -14;
        weight_rom[751] = 4;
        weight_rom[752] = 1;
        weight_rom[753] = -2;
        weight_rom[754] = 2;
        weight_rom[755] = -1;
        weight_rom[756] = 2;
        weight_rom[757] = 1;
        weight_rom[758] = 1;
        weight_rom[759] = -2;
        weight_rom[760] = 0;
        weight_rom[761] = -7;
        weight_rom[762] = -10;
        weight_rom[763] = -6;
        weight_rom[764] = -25;
        weight_rom[765] = -23;
        weight_rom[766] = -27;
        weight_rom[767] = -2;
        weight_rom[768] = -12;
        weight_rom[769] = -33;
        weight_rom[770] = -14;
        weight_rom[771] = -6;
        weight_rom[772] = -12;
        weight_rom[773] = -25;
        weight_rom[774] = -26;
        weight_rom[775] = -20;
        weight_rom[776] = 17;
        weight_rom[777] = 1;
        weight_rom[778] = -2;
        weight_rom[779] = 0;
        weight_rom[780] = -1;
        weight_rom[781] = -2;
        weight_rom[782] = 0;
        weight_rom[783] = 1;
        weight_rom[784] = 0;
        weight_rom[785] = 1;
        weight_rom[786] = 0;
        weight_rom[787] = 0;
        weight_rom[788] = -2;
        weight_rom[789] = 2;
        weight_rom[790] = -1;
        weight_rom[791] = -2;
        weight_rom[792] = 1;
        weight_rom[793] = 1;
        weight_rom[794] = 2;
        weight_rom[795] = 1;
        weight_rom[796] = -2;
        weight_rom[797] = -14;
        weight_rom[798] = -1;
        weight_rom[799] = -1;
        weight_rom[800] = 2;
        weight_rom[801] = 1;
        weight_rom[802] = 0;
        weight_rom[803] = 2;
        weight_rom[804] = -1;
        weight_rom[805] = 1;
        weight_rom[806] = 2;
        weight_rom[807] = 2;
        weight_rom[808] = 0;
        weight_rom[809] = 2;
        weight_rom[810] = -2;
        weight_rom[811] = 1;
        weight_rom[812] = 1;
        weight_rom[813] = 0;
        weight_rom[814] = 0;
        weight_rom[815] = -2;
        weight_rom[816] = -1;
        weight_rom[817] = 0;
        weight_rom[818] = -16;
        weight_rom[819] = -30;
        weight_rom[820] = -26;
        weight_rom[821] = -13;
        weight_rom[822] = -20;
        weight_rom[823] = -28;
        weight_rom[824] = -36;
        weight_rom[825] = -32;
        weight_rom[826] = 1;
        weight_rom[827] = 10;
        weight_rom[828] = -22;
        weight_rom[829] = -3;
        weight_rom[830] = -14;
        weight_rom[831] = -9;
        weight_rom[832] = -7;
        weight_rom[833] = -19;
        weight_rom[834] = -18;
        weight_rom[835] = -12;
        weight_rom[836] = 1;
        weight_rom[837] = -1;
        weight_rom[838] = -2;
        weight_rom[839] = 0;
        weight_rom[840] = -1;
        weight_rom[841] = 0;
        weight_rom[842] = 1;
        weight_rom[843] = -1;
        weight_rom[844] = -14;
        weight_rom[845] = -1;
        weight_rom[846] = -25;
        weight_rom[847] = -46;
        weight_rom[848] = -53;
        weight_rom[849] = -60;
        weight_rom[850] = -85;
        weight_rom[851] = -89;
        weight_rom[852] = -101;
        weight_rom[853] = -96;
        weight_rom[854] = -101;
        weight_rom[855] = -68;
        weight_rom[856] = -69;
        weight_rom[857] = -53;
        weight_rom[858] = -36;
        weight_rom[859] = -2;
        weight_rom[860] = -15;
        weight_rom[861] = -15;
        weight_rom[862] = -4;
        weight_rom[863] = -19;
        weight_rom[864] = -6;
        weight_rom[865] = -12;
        weight_rom[866] = -1;
        weight_rom[867] = 2;
        weight_rom[868] = 0;
        weight_rom[869] = 0;
        weight_rom[870] = 1;
        weight_rom[871] = 2;
        weight_rom[872] = 0;
        weight_rom[873] = -8;
        weight_rom[874] = -20;
        weight_rom[875] = -36;
        weight_rom[876] = -29;
        weight_rom[877] = -23;
        weight_rom[878] = -17;
        weight_rom[879] = -18;
        weight_rom[880] = -20;
        weight_rom[881] = -40;
        weight_rom[882] = -22;
        weight_rom[883] = -32;
        weight_rom[884] = -29;
        weight_rom[885] = -22;
        weight_rom[886] = -16;
        weight_rom[887] = -19;
        weight_rom[888] = -17;
        weight_rom[889] = -1;
        weight_rom[890] = -12;
        weight_rom[891] = -12;
        weight_rom[892] = -42;
        weight_rom[893] = -13;
        weight_rom[894] = 2;
        weight_rom[895] = 0;
        weight_rom[896] = 2;
        weight_rom[897] = 0;
        weight_rom[898] = 0;
        weight_rom[899] = 0;
        weight_rom[900] = 5;
        weight_rom[901] = 7;
        weight_rom[902] = 10;
        weight_rom[903] = 24;
        weight_rom[904] = 10;
        weight_rom[905] = 16;
        weight_rom[906] = 5;
        weight_rom[907] = 19;
        weight_rom[908] = 6;
        weight_rom[909] = 2;
        weight_rom[910] = 3;
        weight_rom[911] = -3;
        weight_rom[912] = 2;
        weight_rom[913] = -1;
        weight_rom[914] = 2;
        weight_rom[915] = 1;
        weight_rom[916] = -1;
        weight_rom[917] = 6;
        weight_rom[918] = -5;
        weight_rom[919] = 12;
        weight_rom[920] = 29;
        weight_rom[921] = 21;
        weight_rom[922] = 13;
        weight_rom[923] = 1;
        weight_rom[924] = 1;
        weight_rom[925] = -1;
        weight_rom[926] = 0;
        weight_rom[927] = 13;
        weight_rom[928] = -6;
        weight_rom[929] = 17;
        weight_rom[930] = 24;
        weight_rom[931] = 12;
        weight_rom[932] = 16;
        weight_rom[933] = 12;
        weight_rom[934] = 11;
        weight_rom[935] = 7;
        weight_rom[936] = 6;
        weight_rom[937] = 2;
        weight_rom[938] = 2;
        weight_rom[939] = -1;
        weight_rom[940] = -2;
        weight_rom[941] = 2;
        weight_rom[942] = -1;
        weight_rom[943] = -2;
        weight_rom[944] = -1;
        weight_rom[945] = -4;
        weight_rom[946] = 1;
        weight_rom[947] = 16;
        weight_rom[948] = 20;
        weight_rom[949] = 28;
        weight_rom[950] = -3;
        weight_rom[951] = -1;
        weight_rom[952] = 1;
        weight_rom[953] = -2;
        weight_rom[954] = 22;
        weight_rom[955] = 22;
        weight_rom[956] = 14;
        weight_rom[957] = 11;
        weight_rom[958] = 15;
        weight_rom[959] = 2;
        weight_rom[960] = 17;
        weight_rom[961] = 14;
        weight_rom[962] = 16;
        weight_rom[963] = 8;
        weight_rom[964] = 0;
        weight_rom[965] = 0;
        weight_rom[966] = 3;
        weight_rom[967] = 3;
        weight_rom[968] = 5;
        weight_rom[969] = 6;
        weight_rom[970] = 0;
        weight_rom[971] = 1;
        weight_rom[972] = 4;
        weight_rom[973] = -4;
        weight_rom[974] = 5;
        weight_rom[975] = 10;
        weight_rom[976] = 24;
        weight_rom[977] = 25;
        weight_rom[978] = 10;
        weight_rom[979] = -27;
        weight_rom[980] = -1;
        weight_rom[981] = -11;
        weight_rom[982] = 6;
        weight_rom[983] = 17;
        weight_rom[984] = 4;
        weight_rom[985] = 8;
        weight_rom[986] = 4;
        weight_rom[987] = 2;
        weight_rom[988] = 4;
        weight_rom[989] = 7;
        weight_rom[990] = 6;
        weight_rom[991] = 1;
        weight_rom[992] = 0;
        weight_rom[993] = 2;
        weight_rom[994] = 2;
        weight_rom[995] = 7;
        weight_rom[996] = 7;
        weight_rom[997] = 6;
        weight_rom[998] = 0;
        weight_rom[999] = 6;
        weight_rom[1000] = 2;
        weight_rom[1001] = 0;
        weight_rom[1002] = 1;
        weight_rom[1003] = 5;
        weight_rom[1004] = 8;
        weight_rom[1005] = 30;
        weight_rom[1006] = 1;
        weight_rom[1007] = -16;
        weight_rom[1008] = 11;
        weight_rom[1009] = 17;
        weight_rom[1010] = 18;
        weight_rom[1011] = 15;
        weight_rom[1012] = 11;
        weight_rom[1013] = 18;
        weight_rom[1014] = 3;
        weight_rom[1015] = 5;
        weight_rom[1016] = 4;
        weight_rom[1017] = 1;
        weight_rom[1018] = 4;
        weight_rom[1019] = 5;
        weight_rom[1020] = 1;
        weight_rom[1021] = 0;
        weight_rom[1022] = -3;
        weight_rom[1023] = -3;
        weight_rom[1024] = 0;
        weight_rom[1025] = -1;
        weight_rom[1026] = 1;
        weight_rom[1027] = 2;
        weight_rom[1028] = 8;
        weight_rom[1029] = 4;
        weight_rom[1030] = 3;
        weight_rom[1031] = 4;
        weight_rom[1032] = 31;
        weight_rom[1033] = 24;
        weight_rom[1034] = 3;
        weight_rom[1035] = -20;
        weight_rom[1036] = 18;
        weight_rom[1037] = 31;
        weight_rom[1038] = 44;
        weight_rom[1039] = 31;
        weight_rom[1040] = 8;
        weight_rom[1041] = 10;
        weight_rom[1042] = 6;
        weight_rom[1043] = -1;
        weight_rom[1044] = -2;
        weight_rom[1045] = 4;
        weight_rom[1046] = 5;
        weight_rom[1047] = 7;
        weight_rom[1048] = 7;
        weight_rom[1049] = -3;
        weight_rom[1050] = -9;
        weight_rom[1051] = 1;
        weight_rom[1052] = 2;
        weight_rom[1053] = 6;
        weight_rom[1054] = 3;
        weight_rom[1055] = 7;
        weight_rom[1056] = 9;
        weight_rom[1057] = 10;
        weight_rom[1058] = 10;
        weight_rom[1059] = -3;
        weight_rom[1060] = 12;
        weight_rom[1061] = 27;
        weight_rom[1062] = 11;
        weight_rom[1063] = 17;
        weight_rom[1064] = 18;
        weight_rom[1065] = 18;
        weight_rom[1066] = 42;
        weight_rom[1067] = 33;
        weight_rom[1068] = 2;
        weight_rom[1069] = -7;
        weight_rom[1070] = -6;
        weight_rom[1071] = 4;
        weight_rom[1072] = 4;
        weight_rom[1073] = 3;
        weight_rom[1074] = 8;
        weight_rom[1075] = 7;
        weight_rom[1076] = 4;
        weight_rom[1077] = -4;
        weight_rom[1078] = -12;
        weight_rom[1079] = -3;
        weight_rom[1080] = 11;
        weight_rom[1081] = 9;
        weight_rom[1082] = 4;
        weight_rom[1083] = 8;
        weight_rom[1084] = 5;
        weight_rom[1085] = 12;
        weight_rom[1086] = 5;
        weight_rom[1087] = -1;
        weight_rom[1088] = 13;
        weight_rom[1089] = 48;
        weight_rom[1090] = 28;
        weight_rom[1091] = 13;
        weight_rom[1092] = 21;
        weight_rom[1093] = 35;
        weight_rom[1094] = 60;
        weight_rom[1095] = 24;
        weight_rom[1096] = 7;
        weight_rom[1097] = 2;
        weight_rom[1098] = 11;
        weight_rom[1099] = 0;
        weight_rom[1100] = 1;
        weight_rom[1101] = 9;
        weight_rom[1102] = 10;
        weight_rom[1103] = 16;
        weight_rom[1104] = 10;
        weight_rom[1105] = 2;
        weight_rom[1106] = -3;
        weight_rom[1107] = 7;
        weight_rom[1108] = 18;
        weight_rom[1109] = 27;
        weight_rom[1110] = 8;
        weight_rom[1111] = 10;
        weight_rom[1112] = 9;
        weight_rom[1113] = 4;
        weight_rom[1114] = 5;
        weight_rom[1115] = -17;
        weight_rom[1116] = -11;
        weight_rom[1117] = 21;
        weight_rom[1118] = 8;
        weight_rom[1119] = -2;
        weight_rom[1120] = 17;
        weight_rom[1121] = 19;
        weight_rom[1122] = 44;
        weight_rom[1123] = 17;
        weight_rom[1124] = 21;
        weight_rom[1125] = 7;
        weight_rom[1126] = 8;
        weight_rom[1127] = 3;
        weight_rom[1128] = 13;
        weight_rom[1129] = 4;
        weight_rom[1130] = 7;
        weight_rom[1131] = 10;
        weight_rom[1132] = 7;
        weight_rom[1133] = 7;
        weight_rom[1134] = -6;
        weight_rom[1135] = 6;
        weight_rom[1136] = 20;
        weight_rom[1137] = 31;
        weight_rom[1138] = 18;
        weight_rom[1139] = 9;
        weight_rom[1140] = 3;
        weight_rom[1141] = -11;
        weight_rom[1142] = -8;
        weight_rom[1143] = -20;
        weight_rom[1144] = -17;
        weight_rom[1145] = 10;
        weight_rom[1146] = 1;
        weight_rom[1147] = -1;
        weight_rom[1148] = -2;
        weight_rom[1149] = -3;
        weight_rom[1150] = 40;
        weight_rom[1151] = 11;
        weight_rom[1152] = 52;
        weight_rom[1153] = 30;
        weight_rom[1154] = 13;
        weight_rom[1155] = 19;
        weight_rom[1156] = 7;
        weight_rom[1157] = 7;
        weight_rom[1158] = 4;
        weight_rom[1159] = 8;
        weight_rom[1160] = 14;
        weight_rom[1161] = 11;
        weight_rom[1162] = -10;
        weight_rom[1163] = 9;
        weight_rom[1164] = 23;
        weight_rom[1165] = 33;
        weight_rom[1166] = 19;
        weight_rom[1167] = 4;
        weight_rom[1168] = 1;
        weight_rom[1169] = -2;
        weight_rom[1170] = -11;
        weight_rom[1171] = -37;
        weight_rom[1172] = -12;
        weight_rom[1173] = -16;
        weight_rom[1174] = -12;
        weight_rom[1175] = -17;
        weight_rom[1176] = 2;
        weight_rom[1177] = 16;
        weight_rom[1178] = 10;
        weight_rom[1179] = 20;
        weight_rom[1180] = 51;
        weight_rom[1181] = 16;
        weight_rom[1182] = 12;
        weight_rom[1183] = 3;
        weight_rom[1184] = 4;
        weight_rom[1185] = 0;
        weight_rom[1186] = -4;
        weight_rom[1187] = -1;
        weight_rom[1188] = 15;
        weight_rom[1189] = 1;
        weight_rom[1190] = 0;
        weight_rom[1191] = 3;
        weight_rom[1192] = 24;
        weight_rom[1193] = 34;
        weight_rom[1194] = 14;
        weight_rom[1195] = 6;
        weight_rom[1196] = 4;
        weight_rom[1197] = -2;
        weight_rom[1198] = -6;
        weight_rom[1199] = -21;
        weight_rom[1200] = -16;
        weight_rom[1201] = -15;
        weight_rom[1202] = -35;
        weight_rom[1203] = -2;
        weight_rom[1204] = 0;
        weight_rom[1205] = -3;
        weight_rom[1206] = 6;
        weight_rom[1207] = 12;
        weight_rom[1208] = 10;
        weight_rom[1209] = -10;
        weight_rom[1210] = 7;
        weight_rom[1211] = 1;
        weight_rom[1212] = -5;
        weight_rom[1213] = -4;
        weight_rom[1214] = -9;
        weight_rom[1215] = 4;
        weight_rom[1216] = 18;
        weight_rom[1217] = -1;
        weight_rom[1218] = -2;
        weight_rom[1219] = 6;
        weight_rom[1220] = 26;
        weight_rom[1221] = 28;
        weight_rom[1222] = 10;
        weight_rom[1223] = -2;
        weight_rom[1224] = 1;
        weight_rom[1225] = 2;
        weight_rom[1226] = 0;
        weight_rom[1227] = -3;
        weight_rom[1228] = -30;
        weight_rom[1229] = -45;
        weight_rom[1230] = 3;
        weight_rom[1231] = -6;
        weight_rom[1232] = 1;
        weight_rom[1233] = 2;
        weight_rom[1234] = 27;
        weight_rom[1235] = 10;
        weight_rom[1236] = -3;
        weight_rom[1237] = -19;
        weight_rom[1238] = -6;
        weight_rom[1239] = -4;
        weight_rom[1240] = 3;
        weight_rom[1241] = -2;
        weight_rom[1242] = -10;
        weight_rom[1243] = 9;
        weight_rom[1244] = 20;
        weight_rom[1245] = 1;
        weight_rom[1246] = -5;
        weight_rom[1247] = 12;
        weight_rom[1248] = 30;
        weight_rom[1249] = 16;
        weight_rom[1250] = 0;
        weight_rom[1251] = -3;
        weight_rom[1252] = -8;
        weight_rom[1253] = -10;
        weight_rom[1254] = -8;
        weight_rom[1255] = -9;
        weight_rom[1256] = -19;
        weight_rom[1257] = -45;
        weight_rom[1258] = -31;
        weight_rom[1259] = 8;
        weight_rom[1260] = 0;
        weight_rom[1261] = 13;
        weight_rom[1262] = 3;
        weight_rom[1263] = 13;
        weight_rom[1264] = -1;
        weight_rom[1265] = -20;
        weight_rom[1266] = -12;
        weight_rom[1267] = -20;
        weight_rom[1268] = -11;
        weight_rom[1269] = -3;
        weight_rom[1270] = -5;
        weight_rom[1271] = 11;
        weight_rom[1272] = 10;
        weight_rom[1273] = 3;
        weight_rom[1274] = 7;
        weight_rom[1275] = 21;
        weight_rom[1276] = 16;
        weight_rom[1277] = 6;
        weight_rom[1278] = -8;
        weight_rom[1279] = -5;
        weight_rom[1280] = -11;
        weight_rom[1281] = 5;
        weight_rom[1282] = -11;
        weight_rom[1283] = 1;
        weight_rom[1284] = -15;
        weight_rom[1285] = -37;
        weight_rom[1286] = -43;
        weight_rom[1287] = -2;
        weight_rom[1288] = 2;
        weight_rom[1289] = 12;
        weight_rom[1290] = 19;
        weight_rom[1291] = 24;
        weight_rom[1292] = -3;
        weight_rom[1293] = -12;
        weight_rom[1294] = 7;
        weight_rom[1295] = -15;
        weight_rom[1296] = -23;
        weight_rom[1297] = -19;
        weight_rom[1298] = -21;
        weight_rom[1299] = -18;
        weight_rom[1300] = -19;
        weight_rom[1301] = -7;
        weight_rom[1302] = -4;
        weight_rom[1303] = 5;
        weight_rom[1304] = -3;
        weight_rom[1305] = -6;
        weight_rom[1306] = -8;
        weight_rom[1307] = -6;
        weight_rom[1308] = -5;
        weight_rom[1309] = -10;
        weight_rom[1310] = -9;
        weight_rom[1311] = -16;
        weight_rom[1312] = -41;
        weight_rom[1313] = -52;
        weight_rom[1314] = -1;
        weight_rom[1315] = -1;
        weight_rom[1316] = -1;
        weight_rom[1317] = 12;
        weight_rom[1318] = 29;
        weight_rom[1319] = 36;
        weight_rom[1320] = 1;
        weight_rom[1321] = 5;
        weight_rom[1322] = 0;
        weight_rom[1323] = -3;
        weight_rom[1324] = -7;
        weight_rom[1325] = -17;
        weight_rom[1326] = -26;
        weight_rom[1327] = -42;
        weight_rom[1328] = -40;
        weight_rom[1329] = -28;
        weight_rom[1330] = -15;
        weight_rom[1331] = -11;
        weight_rom[1332] = -10;
        weight_rom[1333] = -4;
        weight_rom[1334] = -5;
        weight_rom[1335] = 0;
        weight_rom[1336] = -3;
        weight_rom[1337] = -8;
        weight_rom[1338] = -6;
        weight_rom[1339] = -11;
        weight_rom[1340] = -13;
        weight_rom[1341] = -22;
        weight_rom[1342] = -31;
        weight_rom[1343] = -1;
        weight_rom[1344] = 0;
        weight_rom[1345] = 13;
        weight_rom[1346] = 19;
        weight_rom[1347] = 26;
        weight_rom[1348] = 1;
        weight_rom[1349] = 6;
        weight_rom[1350] = 3;
        weight_rom[1351] = -2;
        weight_rom[1352] = -2;
        weight_rom[1353] = -6;
        weight_rom[1354] = -15;
        weight_rom[1355] = -18;
        weight_rom[1356] = -17;
        weight_rom[1357] = -13;
        weight_rom[1358] = -7;
        weight_rom[1359] = -7;
        weight_rom[1360] = -8;
        weight_rom[1361] = 1;
        weight_rom[1362] = -4;
        weight_rom[1363] = 1;
        weight_rom[1364] = -1;
        weight_rom[1365] = -9;
        weight_rom[1366] = -1;
        weight_rom[1367] = -12;
        weight_rom[1368] = -31;
        weight_rom[1369] = 6;
        weight_rom[1370] = -25;
        weight_rom[1371] = -2;
        weight_rom[1372] = 2;
        weight_rom[1373] = 0;
        weight_rom[1374] = 15;
        weight_rom[1375] = 9;
        weight_rom[1376] = 16;
        weight_rom[1377] = 1;
        weight_rom[1378] = 7;
        weight_rom[1379] = -2;
        weight_rom[1380] = -7;
        weight_rom[1381] = -10;
        weight_rom[1382] = -11;
        weight_rom[1383] = -15;
        weight_rom[1384] = -5;
        weight_rom[1385] = -10;
        weight_rom[1386] = -10;
        weight_rom[1387] = -9;
        weight_rom[1388] = -5;
        weight_rom[1389] = -6;
        weight_rom[1390] = -6;
        weight_rom[1391] = -3;
        weight_rom[1392] = -5;
        weight_rom[1393] = -2;
        weight_rom[1394] = -3;
        weight_rom[1395] = -21;
        weight_rom[1396] = -17;
        weight_rom[1397] = -18;
        weight_rom[1398] = -20;
        weight_rom[1399] = 1;
        weight_rom[1400] = 2;
        weight_rom[1401] = -2;
        weight_rom[1402] = 25;
        weight_rom[1403] = 23;
        weight_rom[1404] = 9;
        weight_rom[1405] = 0;
        weight_rom[1406] = -15;
        weight_rom[1407] = -9;
        weight_rom[1408] = -8;
        weight_rom[1409] = -11;
        weight_rom[1410] = -6;
        weight_rom[1411] = 0;
        weight_rom[1412] = 0;
        weight_rom[1413] = -1;
        weight_rom[1414] = -9;
        weight_rom[1415] = -9;
        weight_rom[1416] = -8;
        weight_rom[1417] = -4;
        weight_rom[1418] = -12;
        weight_rom[1419] = -3;
        weight_rom[1420] = -13;
        weight_rom[1421] = -14;
        weight_rom[1422] = -8;
        weight_rom[1423] = -3;
        weight_rom[1424] = -10;
        weight_rom[1425] = -12;
        weight_rom[1426] = -18;
        weight_rom[1427] = 1;
        weight_rom[1428] = 1;
        weight_rom[1429] = -1;
        weight_rom[1430] = -13;
        weight_rom[1431] = 15;
        weight_rom[1432] = 9;
        weight_rom[1433] = -8;
        weight_rom[1434] = -14;
        weight_rom[1435] = -9;
        weight_rom[1436] = -9;
        weight_rom[1437] = -11;
        weight_rom[1438] = -7;
        weight_rom[1439] = -1;
        weight_rom[1440] = -2;
        weight_rom[1441] = -5;
        weight_rom[1442] = -2;
        weight_rom[1443] = -12;
        weight_rom[1444] = -10;
        weight_rom[1445] = -4;
        weight_rom[1446] = -7;
        weight_rom[1447] = -3;
        weight_rom[1448] = -15;
        weight_rom[1449] = -8;
        weight_rom[1450] = -7;
        weight_rom[1451] = 6;
        weight_rom[1452] = 0;
        weight_rom[1453] = -13;
        weight_rom[1454] = -2;
        weight_rom[1455] = -1;
        weight_rom[1456] = -2;
        weight_rom[1457] = 1;
        weight_rom[1458] = -14;
        weight_rom[1459] = 18;
        weight_rom[1460] = 15;
        weight_rom[1461] = 18;
        weight_rom[1462] = 0;
        weight_rom[1463] = 9;
        weight_rom[1464] = 7;
        weight_rom[1465] = -8;
        weight_rom[1466] = 2;
        weight_rom[1467] = 5;
        weight_rom[1468] = -6;
        weight_rom[1469] = -2;
        weight_rom[1470] = -7;
        weight_rom[1471] = -6;
        weight_rom[1472] = -1;
        weight_rom[1473] = 4;
        weight_rom[1474] = 9;
        weight_rom[1475] = 23;
        weight_rom[1476] = 34;
        weight_rom[1477] = 24;
        weight_rom[1478] = 18;
        weight_rom[1479] = 35;
        weight_rom[1480] = 2;
        weight_rom[1481] = -26;
        weight_rom[1482] = -2;
        weight_rom[1483] = -1;
        weight_rom[1484] = 2;
        weight_rom[1485] = -1;
        weight_rom[1486] = 1;
        weight_rom[1487] = -6;
        weight_rom[1488] = 25;
        weight_rom[1489] = 67;
        weight_rom[1490] = 56;
        weight_rom[1491] = 65;
        weight_rom[1492] = 48;
        weight_rom[1493] = 58;
        weight_rom[1494] = 39;
        weight_rom[1495] = 41;
        weight_rom[1496] = 41;
        weight_rom[1497] = 43;
        weight_rom[1498] = 40;
        weight_rom[1499] = 48;
        weight_rom[1500] = 66;
        weight_rom[1501] = 65;
        weight_rom[1502] = 81;
        weight_rom[1503] = 88;
        weight_rom[1504] = 70;
        weight_rom[1505] = 88;
        weight_rom[1506] = 44;
        weight_rom[1507] = 53;
        weight_rom[1508] = 27;
        weight_rom[1509] = -1;
        weight_rom[1510] = -2;
        weight_rom[1511] = 2;
        weight_rom[1512] = -2;
        weight_rom[1513] = -2;
        weight_rom[1514] = 2;
        weight_rom[1515] = 0;
        weight_rom[1516] = 30;
        weight_rom[1517] = 53;
        weight_rom[1518] = 58;
        weight_rom[1519] = 78;
        weight_rom[1520] = 108;
        weight_rom[1521] = 101;
        weight_rom[1522] = 96;
        weight_rom[1523] = 107;
        weight_rom[1524] = 95;
        weight_rom[1525] = 121;
        weight_rom[1526] = 127;
        weight_rom[1527] = 108;
        weight_rom[1528] = 115;
        weight_rom[1529] = 98;
        weight_rom[1530] = 77;
        weight_rom[1531] = 67;
        weight_rom[1532] = 51;
        weight_rom[1533] = 46;
        weight_rom[1534] = 37;
        weight_rom[1535] = 18;
        weight_rom[1536] = -1;
        weight_rom[1537] = -1;
        weight_rom[1538] = 2;
        weight_rom[1539] = -1;
        weight_rom[1540] = -1;
        weight_rom[1541] = 0;
        weight_rom[1542] = 0;
        weight_rom[1543] = 2;
        weight_rom[1544] = -2;
        weight_rom[1545] = 23;
        weight_rom[1546] = 39;
        weight_rom[1547] = 50;
        weight_rom[1548] = 49;
        weight_rom[1549] = 52;
        weight_rom[1550] = 52;
        weight_rom[1551] = 36;
        weight_rom[1552] = 56;
        weight_rom[1553] = 92;
        weight_rom[1554] = 89;
        weight_rom[1555] = 78;
        weight_rom[1556] = 70;
        weight_rom[1557] = 74;
        weight_rom[1558] = 60;
        weight_rom[1559] = 32;
        weight_rom[1560] = 9;
        weight_rom[1561] = 5;
        weight_rom[1562] = 28;
        weight_rom[1563] = 0;
        weight_rom[1564] = 1;
        weight_rom[1565] = 1;
        weight_rom[1566] = -1;
        weight_rom[1567] = 1;
        weight_rom[1568] = -2;
        weight_rom[1569] = -1;
        weight_rom[1570] = -2;
        weight_rom[1571] = -2;
        weight_rom[1572] = 1;
        weight_rom[1573] = 0;
        weight_rom[1574] = -2;
        weight_rom[1575] = 2;
        weight_rom[1576] = 0;
        weight_rom[1577] = 0;
        weight_rom[1578] = 1;
        weight_rom[1579] = 1;
        weight_rom[1580] = -1;
        weight_rom[1581] = 9;
        weight_rom[1582] = 17;
        weight_rom[1583] = 1;
        weight_rom[1584] = -2;
        weight_rom[1585] = 1;
        weight_rom[1586] = 0;
        weight_rom[1587] = 2;
        weight_rom[1588] = -2;
        weight_rom[1589] = -1;
        weight_rom[1590] = 0;
        weight_rom[1591] = 0;
        weight_rom[1592] = 2;
        weight_rom[1593] = -1;
        weight_rom[1594] = 1;
        weight_rom[1595] = 0;
        weight_rom[1596] = 0;
        weight_rom[1597] = 0;
        weight_rom[1598] = 1;
        weight_rom[1599] = 0;
        weight_rom[1600] = 2;
        weight_rom[1601] = -2;
        weight_rom[1602] = -5;
        weight_rom[1603] = -9;
        weight_rom[1604] = -12;
        weight_rom[1605] = -19;
        weight_rom[1606] = -8;
        weight_rom[1607] = -23;
        weight_rom[1608] = -32;
        weight_rom[1609] = -25;
        weight_rom[1610] = 16;
        weight_rom[1611] = 7;
        weight_rom[1612] = 37;
        weight_rom[1613] = 14;
        weight_rom[1614] = -30;
        weight_rom[1615] = 15;
        weight_rom[1616] = 2;
        weight_rom[1617] = -12;
        weight_rom[1618] = -6;
        weight_rom[1619] = 0;
        weight_rom[1620] = 1;
        weight_rom[1621] = -2;
        weight_rom[1622] = 2;
        weight_rom[1623] = 0;
        weight_rom[1624] = -2;
        weight_rom[1625] = 2;
        weight_rom[1626] = -1;
        weight_rom[1627] = 0;
        weight_rom[1628] = -13;
        weight_rom[1629] = 0;
        weight_rom[1630] = -14;
        weight_rom[1631] = -13;
        weight_rom[1632] = 3;
        weight_rom[1633] = 27;
        weight_rom[1634] = -3;
        weight_rom[1635] = 21;
        weight_rom[1636] = 22;
        weight_rom[1637] = 31;
        weight_rom[1638] = 29;
        weight_rom[1639] = 38;
        weight_rom[1640] = 44;
        weight_rom[1641] = 36;
        weight_rom[1642] = 22;
        weight_rom[1643] = 16;
        weight_rom[1644] = 20;
        weight_rom[1645] = 2;
        weight_rom[1646] = -17;
        weight_rom[1647] = 25;
        weight_rom[1648] = 22;
        weight_rom[1649] = 17;
        weight_rom[1650] = 1;
        weight_rom[1651] = 2;
        weight_rom[1652] = -2;
        weight_rom[1653] = 1;
        weight_rom[1654] = -13;
        weight_rom[1655] = -1;
        weight_rom[1656] = 2;
        weight_rom[1657] = 20;
        weight_rom[1658] = -5;
        weight_rom[1659] = 7;
        weight_rom[1660] = 3;
        weight_rom[1661] = 19;
        weight_rom[1662] = 21;
        weight_rom[1663] = 10;
        weight_rom[1664] = 15;
        weight_rom[1665] = 15;
        weight_rom[1666] = 10;
        weight_rom[1667] = 6;
        weight_rom[1668] = 9;
        weight_rom[1669] = 16;
        weight_rom[1670] = 9;
        weight_rom[1671] = 5;
        weight_rom[1672] = 8;
        weight_rom[1673] = -2;
        weight_rom[1674] = -12;
        weight_rom[1675] = -14;
        weight_rom[1676] = -3;
        weight_rom[1677] = 13;
        weight_rom[1678] = 2;
        weight_rom[1679] = 1;
        weight_rom[1680] = 1;
        weight_rom[1681] = 2;
        weight_rom[1682] = 14;
        weight_rom[1683] = -1;
        weight_rom[1684] = -5;
        weight_rom[1685] = 18;
        weight_rom[1686] = 32;
        weight_rom[1687] = 16;
        weight_rom[1688] = 19;
        weight_rom[1689] = 23;
        weight_rom[1690] = 29;
        weight_rom[1691] = 19;
        weight_rom[1692] = 23;
        weight_rom[1693] = 23;
        weight_rom[1694] = 19;
        weight_rom[1695] = 12;
        weight_rom[1696] = 4;
        weight_rom[1697] = 0;
        weight_rom[1698] = 5;
        weight_rom[1699] = -1;
        weight_rom[1700] = 3;
        weight_rom[1701] = -17;
        weight_rom[1702] = -8;
        weight_rom[1703] = -21;
        weight_rom[1704] = -25;
        weight_rom[1705] = 14;
        weight_rom[1706] = 19;
        weight_rom[1707] = -1;
        weight_rom[1708] = -1;
        weight_rom[1709] = -1;
        weight_rom[1710] = 1;
        weight_rom[1711] = 20;
        weight_rom[1712] = 19;
        weight_rom[1713] = 29;
        weight_rom[1714] = 16;
        weight_rom[1715] = 26;
        weight_rom[1716] = 18;
        weight_rom[1717] = 20;
        weight_rom[1718] = 12;
        weight_rom[1719] = 13;
        weight_rom[1720] = 18;
        weight_rom[1721] = 16;
        weight_rom[1722] = 13;
        weight_rom[1723] = 10;
        weight_rom[1724] = 4;
        weight_rom[1725] = -3;
        weight_rom[1726] = -5;
        weight_rom[1727] = -5;
        weight_rom[1728] = -7;
        weight_rom[1729] = -13;
        weight_rom[1730] = -5;
        weight_rom[1731] = -4;
        weight_rom[1732] = -3;
        weight_rom[1733] = 10;
        weight_rom[1734] = 19;
        weight_rom[1735] = -2;
        weight_rom[1736] = -1;
        weight_rom[1737] = 0;
        weight_rom[1738] = -12;
        weight_rom[1739] = 23;
        weight_rom[1740] = 20;
        weight_rom[1741] = 7;
        weight_rom[1742] = 13;
        weight_rom[1743] = 12;
        weight_rom[1744] = 13;
        weight_rom[1745] = 15;
        weight_rom[1746] = 10;
        weight_rom[1747] = 9;
        weight_rom[1748] = 7;
        weight_rom[1749] = 13;
        weight_rom[1750] = 12;
        weight_rom[1751] = 12;
        weight_rom[1752] = 11;
        weight_rom[1753] = 7;
        weight_rom[1754] = 3;
        weight_rom[1755] = -7;
        weight_rom[1756] = -7;
        weight_rom[1757] = -18;
        weight_rom[1758] = -17;
        weight_rom[1759] = -10;
        weight_rom[1760] = -2;
        weight_rom[1761] = 14;
        weight_rom[1762] = 17;
        weight_rom[1763] = 5;
        weight_rom[1764] = 0;
        weight_rom[1765] = 24;
        weight_rom[1766] = 7;
        weight_rom[1767] = 25;
        weight_rom[1768] = 36;
        weight_rom[1769] = 10;
        weight_rom[1770] = 9;
        weight_rom[1771] = -3;
        weight_rom[1772] = 4;
        weight_rom[1773] = -5;
        weight_rom[1774] = -1;
        weight_rom[1775] = -5;
        weight_rom[1776] = -2;
        weight_rom[1777] = 4;
        weight_rom[1778] = 12;
        weight_rom[1779] = 11;
        weight_rom[1780] = 7;
        weight_rom[1781] = -1;
        weight_rom[1782] = -6;
        weight_rom[1783] = -2;
        weight_rom[1784] = 0;
        weight_rom[1785] = -5;
        weight_rom[1786] = -2;
        weight_rom[1787] = -14;
        weight_rom[1788] = -3;
        weight_rom[1789] = 1;
        weight_rom[1790] = 14;
        weight_rom[1791] = 5;
        weight_rom[1792] = -14;
        weight_rom[1793] = 2;
        weight_rom[1794] = 4;
        weight_rom[1795] = 21;
        weight_rom[1796] = 39;
        weight_rom[1797] = 7;
        weight_rom[1798] = 8;
        weight_rom[1799] = 1;
        weight_rom[1800] = -7;
        weight_rom[1801] = -8;
        weight_rom[1802] = 0;
        weight_rom[1803] = -5;
        weight_rom[1804] = 1;
        weight_rom[1805] = 6;
        weight_rom[1806] = 10;
        weight_rom[1807] = 4;
        weight_rom[1808] = -1;
        weight_rom[1809] = -1;
        weight_rom[1810] = -1;
        weight_rom[1811] = 0;
        weight_rom[1812] = 1;
        weight_rom[1813] = 5;
        weight_rom[1814] = 5;
        weight_rom[1815] = -19;
        weight_rom[1816] = -14;
        weight_rom[1817] = 9;
        weight_rom[1818] = 27;
        weight_rom[1819] = 14;
        weight_rom[1820] = 6;
        weight_rom[1821] = 11;
        weight_rom[1822] = -28;
        weight_rom[1823] = 30;
        weight_rom[1824] = 35;
        weight_rom[1825] = 14;
        weight_rom[1826] = 6;
        weight_rom[1827] = -1;
        weight_rom[1828] = -13;
        weight_rom[1829] = -2;
        weight_rom[1830] = -2;
        weight_rom[1831] = -9;
        weight_rom[1832] = -10;
        weight_rom[1833] = -9;
        weight_rom[1834] = -1;
        weight_rom[1835] = 0;
        weight_rom[1836] = -4;
        weight_rom[1837] = 1;
        weight_rom[1838] = 1;
        weight_rom[1839] = 4;
        weight_rom[1840] = 5;
        weight_rom[1841] = 0;
        weight_rom[1842] = 4;
        weight_rom[1843] = -8;
        weight_rom[1844] = -23;
        weight_rom[1845] = -6;
        weight_rom[1846] = 18;
        weight_rom[1847] = 0;
        weight_rom[1848] = 9;
        weight_rom[1849] = 7;
        weight_rom[1850] = -8;
        weight_rom[1851] = 17;
        weight_rom[1852] = 9;
        weight_rom[1853] = 8;
        weight_rom[1854] = 6;
        weight_rom[1855] = 0;
        weight_rom[1856] = -6;
        weight_rom[1857] = -10;
        weight_rom[1858] = -8;
        weight_rom[1859] = -16;
        weight_rom[1860] = -23;
        weight_rom[1861] = -25;
        weight_rom[1862] = -2;
        weight_rom[1863] = 6;
        weight_rom[1864] = 7;
        weight_rom[1865] = 0;
        weight_rom[1866] = 5;
        weight_rom[1867] = 9;
        weight_rom[1868] = 9;
        weight_rom[1869] = 18;
        weight_rom[1870] = 13;
        weight_rom[1871] = -5;
        weight_rom[1872] = -19;
        weight_rom[1873] = -7;
        weight_rom[1874] = 11;
        weight_rom[1875] = 17;
        weight_rom[1876] = 2;
        weight_rom[1877] = 6;
        weight_rom[1878] = -7;
        weight_rom[1879] = 18;
        weight_rom[1880] = 0;
        weight_rom[1881] = -3;
        weight_rom[1882] = -12;
        weight_rom[1883] = -10;
        weight_rom[1884] = -10;
        weight_rom[1885] = -15;
        weight_rom[1886] = -11;
        weight_rom[1887] = -12;
        weight_rom[1888] = -20;
        weight_rom[1889] = -19;
        weight_rom[1890] = 9;
        weight_rom[1891] = 9;
        weight_rom[1892] = 8;
        weight_rom[1893] = 8;
        weight_rom[1894] = 9;
        weight_rom[1895] = 11;
        weight_rom[1896] = 15;
        weight_rom[1897] = 14;
        weight_rom[1898] = 19;
        weight_rom[1899] = -4;
        weight_rom[1900] = 2;
        weight_rom[1901] = -6;
        weight_rom[1902] = -6;
        weight_rom[1903] = 13;
        weight_rom[1904] = -13;
        weight_rom[1905] = -14;
        weight_rom[1906] = -16;
        weight_rom[1907] = -8;
        weight_rom[1908] = -1;
        weight_rom[1909] = -3;
        weight_rom[1910] = -27;
        weight_rom[1911] = -22;
        weight_rom[1912] = -18;
        weight_rom[1913] = -14;
        weight_rom[1914] = -10;
        weight_rom[1915] = -6;
        weight_rom[1916] = -13;
        weight_rom[1917] = -10;
        weight_rom[1918] = 22;
        weight_rom[1919] = 12;
        weight_rom[1920] = 16;
        weight_rom[1921] = 17;
        weight_rom[1922] = 18;
        weight_rom[1923] = 21;
        weight_rom[1924] = 14;
        weight_rom[1925] = 10;
        weight_rom[1926] = -7;
        weight_rom[1927] = -22;
        weight_rom[1928] = -13;
        weight_rom[1929] = 22;
        weight_rom[1930] = 25;
        weight_rom[1931] = 12;
        weight_rom[1932] = 2;
        weight_rom[1933] = -14;
        weight_rom[1934] = -5;
        weight_rom[1935] = -17;
        weight_rom[1936] = -17;
        weight_rom[1937] = -30;
        weight_rom[1938] = -21;
        weight_rom[1939] = -21;
        weight_rom[1940] = -9;
        weight_rom[1941] = -10;
        weight_rom[1942] = -16;
        weight_rom[1943] = -4;
        weight_rom[1944] = -2;
        weight_rom[1945] = 13;
        weight_rom[1946] = 27;
        weight_rom[1947] = 11;
        weight_rom[1948] = 16;
        weight_rom[1949] = 22;
        weight_rom[1950] = 22;
        weight_rom[1951] = 8;
        weight_rom[1952] = -1;
        weight_rom[1953] = -10;
        weight_rom[1954] = -40;
        weight_rom[1955] = -37;
        weight_rom[1956] = -6;
        weight_rom[1957] = 33;
        weight_rom[1958] = 29;
        weight_rom[1959] = -1;
        weight_rom[1960] = -1;
        weight_rom[1961] = 8;
        weight_rom[1962] = -13;
        weight_rom[1963] = -9;
        weight_rom[1964] = -20;
        weight_rom[1965] = -24;
        weight_rom[1966] = -21;
        weight_rom[1967] = -13;
        weight_rom[1968] = -9;
        weight_rom[1969] = -11;
        weight_rom[1970] = -12;
        weight_rom[1971] = 1;
        weight_rom[1972] = 7;
        weight_rom[1973] = 18;
        weight_rom[1974] = 23;
        weight_rom[1975] = 11;
        weight_rom[1976] = 16;
        weight_rom[1977] = 23;
        weight_rom[1978] = 11;
        weight_rom[1979] = -6;
        weight_rom[1980] = -12;
        weight_rom[1981] = -19;
        weight_rom[1982] = -32;
        weight_rom[1983] = -26;
        weight_rom[1984] = -18;
        weight_rom[1985] = 24;
        weight_rom[1986] = 49;
        weight_rom[1987] = 0;
        weight_rom[1988] = 1;
        weight_rom[1989] = 15;
        weight_rom[1990] = -6;
        weight_rom[1991] = 1;
        weight_rom[1992] = 17;
        weight_rom[1993] = -6;
        weight_rom[1994] = -4;
        weight_rom[1995] = -5;
        weight_rom[1996] = -9;
        weight_rom[1997] = -11;
        weight_rom[1998] = -11;
        weight_rom[1999] = 2;
        weight_rom[2000] = 15;
        weight_rom[2001] = 36;
        weight_rom[2002] = 22;
        weight_rom[2003] = 10;
        weight_rom[2004] = 18;
        weight_rom[2005] = 10;
        weight_rom[2006] = -5;
        weight_rom[2007] = -11;
        weight_rom[2008] = -19;
        weight_rom[2009] = -18;
        weight_rom[2010] = -25;
        weight_rom[2011] = -22;
        weight_rom[2012] = 5;
        weight_rom[2013] = 31;
        weight_rom[2014] = 36;
        weight_rom[2015] = 19;
        weight_rom[2016] = -1;
        weight_rom[2017] = -1;
        weight_rom[2018] = 33;
        weight_rom[2019] = 26;
        weight_rom[2020] = 13;
        weight_rom[2021] = 13;
        weight_rom[2022] = 4;
        weight_rom[2023] = 10;
        weight_rom[2024] = -6;
        weight_rom[2025] = 5;
        weight_rom[2026] = 1;
        weight_rom[2027] = 10;
        weight_rom[2028] = 26;
        weight_rom[2029] = 29;
        weight_rom[2030] = 21;
        weight_rom[2031] = 9;
        weight_rom[2032] = 17;
        weight_rom[2033] = 6;
        weight_rom[2034] = -9;
        weight_rom[2035] = -14;
        weight_rom[2036] = -12;
        weight_rom[2037] = -7;
        weight_rom[2038] = -9;
        weight_rom[2039] = 0;
        weight_rom[2040] = 17;
        weight_rom[2041] = 60;
        weight_rom[2042] = 64;
        weight_rom[2043] = 29;
        weight_rom[2044] = -2;
        weight_rom[2045] = 2;
        weight_rom[2046] = 26;
        weight_rom[2047] = 38;
        weight_rom[2048] = 18;
        weight_rom[2049] = 6;
        weight_rom[2050] = -5;
        weight_rom[2051] = -4;
        weight_rom[2052] = -1;
        weight_rom[2053] = 2;
        weight_rom[2054] = 4;
        weight_rom[2055] = 14;
        weight_rom[2056] = 29;
        weight_rom[2057] = 23;
        weight_rom[2058] = 18;
        weight_rom[2059] = 8;
        weight_rom[2060] = 5;
        weight_rom[2061] = -4;
        weight_rom[2062] = -12;
        weight_rom[2063] = -4;
        weight_rom[2064] = -9;
        weight_rom[2065] = 1;
        weight_rom[2066] = 4;
        weight_rom[2067] = 10;
        weight_rom[2068] = 2;
        weight_rom[2069] = 70;
        weight_rom[2070] = 63;
        weight_rom[2071] = 2;
        weight_rom[2072] = 0;
        weight_rom[2073] = 0;
        weight_rom[2074] = 40;
        weight_rom[2075] = 40;
        weight_rom[2076] = 9;
        weight_rom[2077] = 4;
        weight_rom[2078] = -2;
        weight_rom[2079] = -8;
        weight_rom[2080] = -5;
        weight_rom[2081] = -1;
        weight_rom[2082] = 3;
        weight_rom[2083] = 2;
        weight_rom[2084] = 7;
        weight_rom[2085] = 14;
        weight_rom[2086] = 12;
        weight_rom[2087] = 8;
        weight_rom[2088] = 10;
        weight_rom[2089] = 6;
        weight_rom[2090] = 8;
        weight_rom[2091] = 3;
        weight_rom[2092] = 8;
        weight_rom[2093] = 5;
        weight_rom[2094] = 12;
        weight_rom[2095] = 15;
        weight_rom[2096] = 28;
        weight_rom[2097] = 76;
        weight_rom[2098] = 33;
        weight_rom[2099] = 28;
        weight_rom[2100] = 1;
        weight_rom[2101] = 1;
        weight_rom[2102] = 9;
        weight_rom[2103] = 44;
        weight_rom[2104] = 10;
        weight_rom[2105] = 5;
        weight_rom[2106] = 0;
        weight_rom[2107] = 8;
        weight_rom[2108] = -4;
        weight_rom[2109] = 3;
        weight_rom[2110] = -7;
        weight_rom[2111] = -16;
        weight_rom[2112] = -14;
        weight_rom[2113] = -1;
        weight_rom[2114] = 2;
        weight_rom[2115] = 7;
        weight_rom[2116] = 8;
        weight_rom[2117] = 9;
        weight_rom[2118] = 9;
        weight_rom[2119] = 10;
        weight_rom[2120] = 8;
        weight_rom[2121] = 10;
        weight_rom[2122] = 14;
        weight_rom[2123] = 14;
        weight_rom[2124] = 12;
        weight_rom[2125] = 56;
        weight_rom[2126] = 50;
        weight_rom[2127] = 15;
        weight_rom[2128] = 1;
        weight_rom[2129] = -7;
        weight_rom[2130] = 14;
        weight_rom[2131] = 55;
        weight_rom[2132] = 37;
        weight_rom[2133] = 6;
        weight_rom[2134] = 12;
        weight_rom[2135] = 9;
        weight_rom[2136] = 4;
        weight_rom[2137] = 4;
        weight_rom[2138] = -4;
        weight_rom[2139] = -12;
        weight_rom[2140] = -17;
        weight_rom[2141] = -13;
        weight_rom[2142] = -4;
        weight_rom[2143] = 1;
        weight_rom[2144] = 6;
        weight_rom[2145] = 9;
        weight_rom[2146] = 14;
        weight_rom[2147] = 12;
        weight_rom[2148] = 16;
        weight_rom[2149] = 10;
        weight_rom[2150] = 0;
        weight_rom[2151] = 16;
        weight_rom[2152] = 38;
        weight_rom[2153] = 35;
        weight_rom[2154] = 26;
        weight_rom[2155] = 0;
        weight_rom[2156] = 1;
        weight_rom[2157] = 12;
        weight_rom[2158] = 36;
        weight_rom[2159] = 57;
        weight_rom[2160] = 23;
        weight_rom[2161] = 14;
        weight_rom[2162] = 6;
        weight_rom[2163] = 4;
        weight_rom[2164] = 3;
        weight_rom[2165] = -6;
        weight_rom[2166] = -6;
        weight_rom[2167] = -11;
        weight_rom[2168] = -14;
        weight_rom[2169] = -10;
        weight_rom[2170] = -8;
        weight_rom[2171] = -11;
        weight_rom[2172] = -3;
        weight_rom[2173] = 0;
        weight_rom[2174] = 11;
        weight_rom[2175] = 11;
        weight_rom[2176] = 6;
        weight_rom[2177] = 2;
        weight_rom[2178] = 5;
        weight_rom[2179] = 17;
        weight_rom[2180] = 38;
        weight_rom[2181] = 30;
        weight_rom[2182] = 14;
        weight_rom[2183] = 0;
        weight_rom[2184] = 1;
        weight_rom[2185] = 0;
        weight_rom[2186] = 42;
        weight_rom[2187] = 52;
        weight_rom[2188] = 27;
        weight_rom[2189] = 13;
        weight_rom[2190] = 13;
        weight_rom[2191] = 9;
        weight_rom[2192] = -2;
        weight_rom[2193] = -4;
        weight_rom[2194] = -4;
        weight_rom[2195] = 1;
        weight_rom[2196] = -5;
        weight_rom[2197] = -8;
        weight_rom[2198] = -8;
        weight_rom[2199] = -6;
        weight_rom[2200] = -8;
        weight_rom[2201] = 2;
        weight_rom[2202] = -2;
        weight_rom[2203] = 5;
        weight_rom[2204] = 6;
        weight_rom[2205] = 4;
        weight_rom[2206] = 3;
        weight_rom[2207] = 17;
        weight_rom[2208] = 26;
        weight_rom[2209] = 7;
        weight_rom[2210] = 19;
        weight_rom[2211] = 2;
        weight_rom[2212] = 1;
        weight_rom[2213] = 2;
        weight_rom[2214] = 35;
        weight_rom[2215] = 44;
        weight_rom[2216] = 31;
        weight_rom[2217] = 5;
        weight_rom[2218] = 5;
        weight_rom[2219] = -1;
        weight_rom[2220] = 3;
        weight_rom[2221] = 2;
        weight_rom[2222] = -3;
        weight_rom[2223] = 0;
        weight_rom[2224] = 5;
        weight_rom[2225] = 6;
        weight_rom[2226] = -4;
        weight_rom[2227] = -7;
        weight_rom[2228] = -6;
        weight_rom[2229] = -14;
        weight_rom[2230] = 3;
        weight_rom[2231] = 6;
        weight_rom[2232] = 3;
        weight_rom[2233] = 6;
        weight_rom[2234] = 22;
        weight_rom[2235] = 14;
        weight_rom[2236] = 1;
        weight_rom[2237] = -3;
        weight_rom[2238] = 15;
        weight_rom[2239] = 0;
        weight_rom[2240] = -2;
        weight_rom[2241] = -2;
        weight_rom[2242] = 21;
        weight_rom[2243] = 9;
        weight_rom[2244] = 20;
        weight_rom[2245] = 15;
        weight_rom[2246] = 9;
        weight_rom[2247] = 2;
        weight_rom[2248] = 4;
        weight_rom[2249] = 1;
        weight_rom[2250] = 6;
        weight_rom[2251] = 7;
        weight_rom[2252] = 6;
        weight_rom[2253] = 3;
        weight_rom[2254] = 5;
        weight_rom[2255] = 6;
        weight_rom[2256] = 9;
        weight_rom[2257] = 7;
        weight_rom[2258] = 15;
        weight_rom[2259] = 13;
        weight_rom[2260] = 8;
        weight_rom[2261] = 24;
        weight_rom[2262] = 8;
        weight_rom[2263] = 10;
        weight_rom[2264] = 26;
        weight_rom[2265] = 19;
        weight_rom[2266] = 2;
        weight_rom[2267] = -2;
        weight_rom[2268] = -2;
        weight_rom[2269] = -2;
        weight_rom[2270] = 0;
        weight_rom[2271] = -11;
        weight_rom[2272] = -27;
        weight_rom[2273] = -29;
        weight_rom[2274] = -7;
        weight_rom[2275] = -22;
        weight_rom[2276] = 2;
        weight_rom[2277] = 2;
        weight_rom[2278] = 10;
        weight_rom[2279] = 6;
        weight_rom[2280] = 13;
        weight_rom[2281] = 13;
        weight_rom[2282] = 20;
        weight_rom[2283] = 12;
        weight_rom[2284] = 26;
        weight_rom[2285] = 32;
        weight_rom[2286] = 33;
        weight_rom[2287] = 39;
        weight_rom[2288] = 46;
        weight_rom[2289] = 26;
        weight_rom[2290] = -4;
        weight_rom[2291] = 14;
        weight_rom[2292] = 12;
        weight_rom[2293] = 1;
        weight_rom[2294] = -1;
        weight_rom[2295] = -1;
        weight_rom[2296] = -1;
        weight_rom[2297] = 0;
        weight_rom[2298] = -1;
        weight_rom[2299] = 0;
        weight_rom[2300] = -14;
        weight_rom[2301] = -28;
        weight_rom[2302] = -7;
        weight_rom[2303] = -5;
        weight_rom[2304] = 13;
        weight_rom[2305] = 16;
        weight_rom[2306] = -3;
        weight_rom[2307] = -2;
        weight_rom[2308] = 1;
        weight_rom[2309] = 9;
        weight_rom[2310] = 13;
        weight_rom[2311] = 3;
        weight_rom[2312] = 28;
        weight_rom[2313] = 34;
        weight_rom[2314] = 34;
        weight_rom[2315] = 28;
        weight_rom[2316] = 44;
        weight_rom[2317] = 21;
        weight_rom[2318] = 12;
        weight_rom[2319] = 13;
        weight_rom[2320] = -1;
        weight_rom[2321] = -1;
        weight_rom[2322] = 0;
        weight_rom[2323] = 0;
        weight_rom[2324] = 1;
        weight_rom[2325] = -1;
        weight_rom[2326] = -1;
        weight_rom[2327] = 0;
        weight_rom[2328] = 0;
        weight_rom[2329] = -11;
        weight_rom[2330] = 3;
        weight_rom[2331] = 21;
        weight_rom[2332] = 29;
        weight_rom[2333] = 27;
        weight_rom[2334] = 3;
        weight_rom[2335] = 12;
        weight_rom[2336] = 25;
        weight_rom[2337] = 24;
        weight_rom[2338] = 29;
        weight_rom[2339] = 23;
        weight_rom[2340] = 15;
        weight_rom[2341] = 15;
        weight_rom[2342] = 9;
        weight_rom[2343] = 17;
        weight_rom[2344] = -8;
        weight_rom[2345] = -11;
        weight_rom[2346] = -8;
        weight_rom[2347] = -1;
        weight_rom[2348] = -2;
        weight_rom[2349] = -1;
        weight_rom[2350] = -2;
        weight_rom[2351] = 0;
        weight_rom[2352] = 21;
        weight_rom[2353] = 127;
        weight_rom[2354] = -17;
        weight_rom[2355] = -32;
        weight_rom[2356] = -61;
        weight_rom[2357] = -83;
        weight_rom[2358] = -69;
        weight_rom[2359] = -86;
        weight_rom[2360] = 71;
        weight_rom[2361] = 13;
        weight_rom[2362] = -94;
        weight_rom[2363] = 70;
        weight_rom[2364] = -76;
        weight_rom[2365] = 17;
        weight_rom[2366] = 50;
        weight_rom[2367] = 71;
        weight_rom[2368] = 29;
        weight_rom[2369] = -72;
        weight_rom[2370] = 10;
        weight_rom[2371] = 9;
        weight_rom[2372] = -66;
        weight_rom[2373] = 97;
        weight_rom[2374] = -127;
        weight_rom[2375] = -40;
        weight_rom[2376] = -106;
        weight_rom[2377] = 68;
        weight_rom[2378] = 1;
        weight_rom[2379] = 24;
        weight_rom[2380] = -21;
        weight_rom[2381] = 21;
        weight_rom[2382] = -9;
        weight_rom[2383] = 57;
        weight_rom[2384] = -16;
        weight_rom[2385] = 127;
        weight_rom[2386] = 27;
        weight_rom[2387] = -35;
        weight_rom[2388] = -12;
        weight_rom[2389] = -68;
        weight_rom[2390] = 65;
        weight_rom[2391] = -19;
        weight_rom[2392] = -34;
        weight_rom[2393] = -9;
        weight_rom[2394] = -65;
    end

    // 主状态机和MAC单元
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            valid <= 0;
            digit_out <= 0;
            neuron_idx <= 0;
            input_idx <= 0;
            accumulator <= 0;
            layer1_done <= 0;
        end else begin
            case (state)
                IDLE: begin
                    valid <= 0;
                    if (start) begin
                        state <= LAYER1;
                        neuron_idx <= 0;
                        input_idx <= 0;
                        layer1_done <= 0;
                        accumulator <= $signed({{16{weight_rom[2352][7]}}, weight_rom[2352]});
                    end
                end

                LAYER1: begin
                    // Layer1 MAC: acc += weight * input
                    if (input_idx < 784) begin
                        accumulator <= accumulator + ($signed({{16{weight_rom[neuron_idx * 784 + input_idx][7]}}, weight_rom[neuron_idx * 784 + input_idx]}) * $signed({23'b0, image_in[input_idx]}));
                        input_idx <= input_idx + 1;
                    end else begin
                        // ReLU并存储
                        layer1_out[neuron_idx] <= (accumulator[23] == 1'b1) ? 24'b0 : accumulator;

                        if (neuron_idx == 2) begin
                            // Layer1完成
                            state <= LAYER2;
                            neuron_idx <= 0;
                            input_idx <= 0;
                            accumulator <= $signed({{16{weight_rom[2385][7]}}, weight_rom[2385]});
                        end else begin
                            // 下一个神经元
                            neuron_idx <= neuron_idx + 1;
                            input_idx <= 0;
                            accumulator <= $signed({{16{weight_rom[2352 + neuron_idx + 1][7]}}, weight_rom[2352 + neuron_idx + 1]});
                        end
                    end
                end

                LAYER2: begin
                    // Layer2 MAC: acc += (weight * layer1_out) >> 7
                    if (input_idx < 3) begin
                        accumulator <= accumulator + (($signed({{16{weight_rom[2355 + neuron_idx * 3 + input_idx][7]}}, weight_rom[2355 + neuron_idx * 3 + input_idx]}) * layer1_out[input_idx]) >>> 7);
                        input_idx <= input_idx + 1;
                    end else begin
                        // 存储输出
                        layer2_out[neuron_idx] <= accumulator;

                        if (neuron_idx == 9) begin
                            // Layer2完成，进入argmax
                            state <= ARGMAX;
                            neuron_idx <= 0;
                            input_idx <= 0;
                            max_idx <= 0;
                            max_val <= layer2_out[0];
                        end else begin
                            // 下一个神经元
                            neuron_idx <= neuron_idx + 1;
                            input_idx <= 0;
                            accumulator <= $signed({{16{weight_rom[2385 + neuron_idx + 1][7]}}, weight_rom[2385 + neuron_idx + 1]});
                        end
                    end
                end

                ARGMAX: begin
                    // 串行比较查找最大值
                    if (input_idx == 0) begin
                        // 初始化已在LAYER2完成
                        input_idx <= 1;
                    end else if (input_idx < 10) begin
                        if (layer2_out[input_idx] > max_val) begin
                            max_val <= layer2_out[input_idx];
                            max_idx <= input_idx[3:0];
                        end
                        input_idx <= input_idx + 1;
                    end else begin
                        // 完成
                        digit_out <= max_idx;
                        valid <= 1;
                        state <= IDLE;
                        input_idx <= 0;
                    end
                end

                default: state <= IDLE;
            endcase
        end
    end

endmodule
