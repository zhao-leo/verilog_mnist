// MNIST模型测试文件 - 使用真实MNIST数据

`timescale 1ns / 1ps

module mnist_model_test;

    reg clk;
    reg rst;
    reg [783:0] image_in;
    reg start;
    wire [3:0] digit_out;
    wire valid;

    // 实例化模块
    mnist_model uut (
        .clk(clk),
        .rst(rst),
        .image_in(image_in),
        .start(start),
        .digit_out(digit_out),
        .valid(valid)
    );

    // 时钟生成
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // 测试流程
    initial begin
        // 初始化
        rst = 1;
        start = 0;
        image_in = 784'b0;

        #20 rst = 0;

        // 测试用例1: 真实MNIST样本 (标签=7, 期望输出=7)
        #50;
        image_in = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001111111111110000000000000000011111111111111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            start = 1;
            #10 start = 0;

            wait(valid);
            $display("Test 1: Layer1[0]=%d, Layer1[1]=%d, Layer1[2]=%d, Layer1[3]=%d",
                     uut.layer1_out[0], uut.layer1_out[1], uut.layer1_out[2], uut.layer1_out[3]);
            $display("         Layer2[0]=%d, [1]=%d, [2]=%d, [3]=%d, [4]=%d",
                     uut.layer2_out[0], uut.layer2_out[1], uut.layer2_out[2], uut.layer2_out[3], uut.layer2_out[4]);
            $display("         Layer2[5]=%d, [6]=%d, [7]=%d, [8]=%d, [9]=%d",
                     uut.layer2_out[5], uut.layer2_out[6], uut.layer2_out[7], uut.layer2_out[8], uut.layer2_out[9]);
            if (digit_out == 7)
                $display("Test 1 PASSED: Label=7, Expected=7, Got=%d", digit_out);
            else
                $display("Test 1 FAILED: Label=7, Expected=7, Got=%d", digit_out);
    
        // 测试用例2: 真实MNIST样本 (标签=2, 期望输出=2)
        #50;
        image_in = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111100000000001111111111111111110000000000111100000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000011000000000000000000111000011100000000000000000001111111110000000000000000000111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            start = 1;
            #10 start = 0;

            wait(valid);
            $display("Test 2: Layer1[0]=%d, Layer1[1]=%d, Layer1[2]=%d, Layer1[3]=%d",
                     uut.layer1_out[0], uut.layer1_out[1], uut.layer1_out[2], uut.layer1_out[3]);
            $display("         Layer2[0]=%d, [1]=%d, [2]=%d, [3]=%d, [4]=%d",
                     uut.layer2_out[0], uut.layer2_out[1], uut.layer2_out[2], uut.layer2_out[3], uut.layer2_out[4]);
            $display("         Layer2[5]=%d, [6]=%d, [7]=%d, [8]=%d, [9]=%d",
                     uut.layer2_out[5], uut.layer2_out[6], uut.layer2_out[7], uut.layer2_out[8], uut.layer2_out[9]);
            if (digit_out == 2)
                $display("Test 2 PASSED: Label=2, Expected=2, Got=%d", digit_out);
            else
                $display("Test 2 FAILED: Label=2, Expected=2, Got=%d", digit_out);
    
        // 测试用例3: 真实MNIST样本 (标签=1, 期望输出=1)
        #50;
        image_in = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            start = 1;
            #10 start = 0;

            wait(valid);
            $display("Test 3: Layer1[0]=%d, Layer1[1]=%d, Layer1[2]=%d, Layer1[3]=%d",
                     uut.layer1_out[0], uut.layer1_out[1], uut.layer1_out[2], uut.layer1_out[3]);
            $display("         Layer2[0]=%d, [1]=%d, [2]=%d, [3]=%d, [4]=%d",
                     uut.layer2_out[0], uut.layer2_out[1], uut.layer2_out[2], uut.layer2_out[3], uut.layer2_out[4]);
            $display("         Layer2[5]=%d, [6]=%d, [7]=%d, [8]=%d, [9]=%d",
                     uut.layer2_out[5], uut.layer2_out[6], uut.layer2_out[7], uut.layer2_out[8], uut.layer2_out[9]);
            if (digit_out == 1)
                $display("Test 3 PASSED: Label=1, Expected=1, Got=%d", digit_out);
            else
                $display("Test 3 FAILED: Label=1, Expected=1, Got=%d", digit_out);
    
        // 测试用例4: 真实MNIST样本 (标签=0, 期望输出=0)
        #50;
        image_in = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011111110000000000000000000111111111100000000000000001111111111110000000000000000111111110011100000000000000111111000001110000000000000011111000000111000000000000011110000000011100000000000001110000000001110000000000001111000000000110000000000000011100000000111000000000000001110000000111100000000000000011100001111110000000000000000111001111110000000000000000011111111111000000000000000000111111111000000000000000000000111111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            start = 1;
            #10 start = 0;

            wait(valid);
            $display("Test 4: Layer1[0]=%d, Layer1[1]=%d, Layer1[2]=%d, Layer1[3]=%d",
                     uut.layer1_out[0], uut.layer1_out[1], uut.layer1_out[2], uut.layer1_out[3]);
            $display("         Layer2[0]=%d, [1]=%d, [2]=%d, [3]=%d, [4]=%d",
                     uut.layer2_out[0], uut.layer2_out[1], uut.layer2_out[2], uut.layer2_out[3], uut.layer2_out[4]);
            $display("         Layer2[5]=%d, [6]=%d, [7]=%d, [8]=%d, [9]=%d",
                     uut.layer2_out[5], uut.layer2_out[6], uut.layer2_out[7], uut.layer2_out[8], uut.layer2_out[9]);
            if (digit_out == 0)
                $display("Test 4 PASSED: Label=0, Expected=0, Got=%d", digit_out);
            else
                $display("Test 4 FAILED: Label=0, Expected=0, Got=%d", digit_out);
    
        // 测试用例5: 真实MNIST样本 (标签=4, 期望输出=4)
        #50;
        image_in = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000111111111110000000000000000011111000011100000000000000001100000000110000000000000001110000000011000000000000000111000000001100000000000000011000000000110000000000000011100000000110000000000000001100000000011000000000000000110000000011000000000000000010000000011000000000000000001000000001100000000000000000110000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            start = 1;
            #10 start = 0;

            wait(valid);
            $display("Test 5: Layer1[0]=%d, Layer1[1]=%d, Layer1[2]=%d, Layer1[3]=%d",
                     uut.layer1_out[0], uut.layer1_out[1], uut.layer1_out[2], uut.layer1_out[3]);
            $display("         Layer2[0]=%d, [1]=%d, [2]=%d, [3]=%d, [4]=%d",
                     uut.layer2_out[0], uut.layer2_out[1], uut.layer2_out[2], uut.layer2_out[3], uut.layer2_out[4]);
            $display("         Layer2[5]=%d, [6]=%d, [7]=%d, [8]=%d, [9]=%d",
                     uut.layer2_out[5], uut.layer2_out[6], uut.layer2_out[7], uut.layer2_out[8], uut.layer2_out[9]);
            if (digit_out == 4)
                $display("Test 5 PASSED: Label=4, Expected=4, Got=%d", digit_out);
            else
                $display("Test 5 FAILED: Label=4, Expected=4, Got=%d", digit_out);
    
        #100;
        $display("\n所有测试完成");
        $finish;
    end

    // 监控输出
    initial begin
        $monitor("Time=%0t rst=%b start=%b valid=%b digit_out=%d",
                 $time, rst, start, valid, digit_out);
    end

endmodule
