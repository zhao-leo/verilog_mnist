// Handwriting模块测试文件
// 正确模拟ARM控制时钟的开始和停止

`timescale 1ns / 1ps

module handwriting_test;

    reg clk;
    reg rst;
    reg data_in;
    wire busy;
    wire [3:0] digit_out;
    wire result_valid;

    // 用于对比测试的直接mnist_model实例
    reg [783:0] direct_image;
    reg direct_start;
    wire [3:0] direct_digit_out;
    wire direct_valid;

    mnist_model direct_mnist (
        .clk(clk),
        .rst(rst),
        .image_in(direct_image),
        .start(direct_start),
        .digit_out(direct_digit_out),
        .valid(direct_valid)
    );

    // 实例化handwriting模块
    handwriting uut (
        .clk(clk),
        .rst(rst),
        .data_in(data_in),
        .busy(busy),
        .digit_out(digit_out),
        .result_valid(result_valid)
    );

    // 测试图像数据（从mnist_model_test.v复制）
    reg [783:0] test_images [0:4];
    integer expected_results [0:4];
    integer i, test_num;
    integer nonzero_ram, nonzero_expected, j;

    // 初始化测试数据（使用mnist_model_test.v中的真实MNIST样本）
    initial begin
        // 测试用例1: 标签=7
        test_images[0] = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001111111111110000000000000000011111111111111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        expected_results[0] = 7;

        // 测试用例2: 标签=2
        test_images[1] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111100000000001111111111111111110000000000111100000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000011000000000000000000111000011100000000000000000001111111110000000000000000000111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        expected_results[1] = 2;

        // 测试用例3: 标签=1
        test_images[2] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        expected_results[2] = 1;

        // 测试用例4: 标签=0
        test_images[3] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011111110000000000000000000111111111100000000000000001111111111110000000000000000111111110011100000000000000111111000001110000000000000011111000000111000000000000011110000000011100000000000001110000000001110000000000001111000000000110000000000000011100000000111000000000000001110000000111100000000000000011100001111110000000000000000111001111110000000000000000011111111111000000000000000000111111111000000000000000000000111111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        expected_results[3] = 0;

        // 测试用例5: 标签=4
        test_images[4] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000111111111110000000000000000011111000011100000000000000001100000000110000000000000001110000000011000000000000000111000000001100000000000000011000000000110000000000000011100000000110000000000000001100000000011000000000000000110000000011000000000000000010000000011000000000000000001000000001100000000000000000110000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        expected_results[4] = 4;
    end

    // 直接测试mnist_model的任务
    task direct_test;
        input [783:0] image_data;
        input integer expected;
        input integer test_id;
        begin
            // 设置图像数据
            direct_image = image_data;
            direct_start = 1;
            #10 clk = 1;
            #10 clk = 0;
            direct_start = 0;

            // 等待计算完成
            while (direct_valid == 0) begin
                #10 clk = 1;
                #10 clk = 0;
            end

            $display("直接测试%0d: 识别结果=%0d (期望=%0d) %s",
                     test_id, direct_digit_out, expected,
                     (direct_digit_out == expected) ? "PASS" : "FAIL");
        end
    endtask

    // ARM模拟：控制时钟的任务
    task arm_send_data;
        input [783:0] image_data;
        input integer expected;
        input integer test_id;
        begin

            // ARM开始提供时钟并发送数据
            // 关键时序：先设置数据，让数据稳定，然后产生时钟上升沿采样
            for (i = 0; i < 784; i = i + 1) begin
                // 1. 确保时钟为低
                clk = 0;
                #5;  // 等待时钟稳定在低电平

                // 2. 在时钟低电平期间设置数据
                data_in = image_data[i];
                #5;  // 给数据足够的建立时间(setup time)

                // 3. 产生上升沿，FPGA在此采样稳定的数据
                clk = 1;
                #10; // 保持高电平
            end

            // 继续提供时钟等待计算完成
            while (busy == 1) begin
                clk = 0;
                #10;
                clk = 1;
                #10;
            end

            // 计算完成，读取结果
            if (result_valid == 1) begin
                if (digit_out == expected)
                    $display("handwriting测试%0d PASSED: 识别结果=%0d", test_id, digit_out);
                else
                    $display("handwriting测试%0d FAILED: 识别结果=%0d, 期望=%0d", test_id, digit_out, expected);
            end else begin
                $display("handwriting测试%0d ERROR: result_valid=0", test_id);
            end

            // ARM停止时钟
            clk = 0;
            #100; // 停止时钟一段时间
        end
    endtask

    // 测试流程
    initial begin
        // 导出波形文件
        $dumpfile("handwriting_test.vcd");
        $dumpvars(0, handwriting_test);
        
        // 初始化
        clk = 0;
        rst = 0;
        data_in = 0;
        direct_image = 784'b0;
        direct_start = 0;

        $display("=== 先用直接mnist_model测试所有样本 ===");
        for (test_num = 0; test_num < 5; test_num = test_num + 1) begin
            rst = 1;
            #20 rst = 0;
            #20;
            direct_test(test_images[test_num], expected_results[test_num], test_num + 1);
        end

        $display("\n=== 再用handwriting模块测试所有样本 ===");
        // 测试5个样本
        for (test_num = 0; test_num < 5; test_num = test_num + 1) begin
            // 复位
            rst = 1;
            data_in = 0;
            clk = 0;
            #20 rst = 0;
            #40;  // 复位后等待更长时间让状态稳定

            // ARM发送数据
            arm_send_data(test_images[test_num], expected_results[test_num], test_num + 1);
        end

        $display("\n所有测试完成");
        $finish;
    end
endmodule
