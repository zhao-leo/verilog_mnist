// MNIST手写数字识别模型 - Int8量化版本（串行计算架构）
// 架构优化：使用单个MAC单元串行计算，大幅减少逻辑门数量
// 网络结构: 784 → 6 → 10 (隐藏层神经元: 6)
// 输入: 28x28二值图像 (784位)
// 输出: 预测数字 (0-9)
// 时钟周期: ~4780 cycles
// ROM大小: 4780 bytes (Layer1: 4710, Layer2: 70)

module mnist_model(
    input wire clk,
    input wire rst,
    input wire [783:0] image_in,  // 28*28 = 784位输入
    input wire start,
    output reg [3:0] digit_out,   // 输出数字 0-9
    output reg valid
);

    // 状态机
    localparam IDLE = 3'd0;
    localparam LAYER1_COMPUTE = 3'd1;
    localparam LAYER1_ACTIVATE = 3'd2;
    localparam LAYER2_COMPUTE = 3'd3;
    localparam ARGMAX = 3'd4;
    localparam DONE = 3'd5;

    reg [2:0] state;
    reg [4:0] neuron_idx;       // 当前神经元索引
    reg [9:0] input_idx;        // 当前输入索引 (0-783 for layer1)

    // MAC单元
    reg signed [31:0] accumulator; // 累加器（32位，保证数值稳定性）

    // 层输出存储
    reg signed [31:0] layer1_out [0:5];
    reg signed [31:0] layer2_out [0:9];

    // ROM: 存储所有权重和偏置 (4780个Int8参数)
    // synthesis attribute: 强制使用Block RAM而不是分布式RAM
    (* ram_style = "block" *) reg signed [7:0] weight_rom [0:4779];

    // 初始化ROM
    initial begin
        weight_rom[0] = 1;
        weight_rom[1] = 0;
        weight_rom[2] = -3;
        weight_rom[3] = 0;
        weight_rom[4] = 1;
        weight_rom[5] = 0;
        weight_rom[6] = -1;
        weight_rom[7] = 1;
        weight_rom[8] = -2;
        weight_rom[9] = 3;
        weight_rom[10] = -1;
        weight_rom[11] = -2;
        weight_rom[12] = -2;
        weight_rom[13] = 18;
        weight_rom[14] = 22;
        weight_rom[15] = 1;
        weight_rom[16] = 1;
        weight_rom[17] = -3;
        weight_rom[18] = -3;
        weight_rom[19] = 1;
        weight_rom[20] = 2;
        weight_rom[21] = 3;
        weight_rom[22] = -1;
        weight_rom[23] = 0;
        weight_rom[24] = -3;
        weight_rom[25] = -1;
        weight_rom[26] = -2;
        weight_rom[27] = 0;
        weight_rom[28] = 2;
        weight_rom[29] = 1;
        weight_rom[30] = -1;
        weight_rom[31] = 0;
        weight_rom[32] = 3;
        weight_rom[33] = -3;
        weight_rom[34] = 2;
        weight_rom[35] = -1;
        weight_rom[36] = -21;
        weight_rom[37] = -8;
        weight_rom[38] = 26;
        weight_rom[39] = -17;
        weight_rom[40] = -3;
        weight_rom[41] = -22;
        weight_rom[42] = 12;
        weight_rom[43] = 27;
        weight_rom[44] = 54;
        weight_rom[45] = 7;
        weight_rom[46] = -31;
        weight_rom[47] = 21;
        weight_rom[48] = 19;
        weight_rom[49] = 19;
        weight_rom[50] = 31;
        weight_rom[51] = 14;
        weight_rom[52] = -1;
        weight_rom[53] = -2;
        weight_rom[54] = 2;
        weight_rom[55] = -2;
        weight_rom[56] = 3;
        weight_rom[57] = 0;
        weight_rom[58] = 2;
        weight_rom[59] = -3;
        weight_rom[60] = -23;
        weight_rom[61] = 0;
        weight_rom[62] = -5;
        weight_rom[63] = -4;
        weight_rom[64] = -6;
        weight_rom[65] = 25;
        weight_rom[66] = 10;
        weight_rom[67] = 22;
        weight_rom[68] = 30;
        weight_rom[69] = 52;
        weight_rom[70] = 33;
        weight_rom[71] = 39;
        weight_rom[72] = 46;
        weight_rom[73] = 32;
        weight_rom[74] = 2;
        weight_rom[75] = -10;
        weight_rom[76] = -28;
        weight_rom[77] = 9;
        weight_rom[78] = 4;
        weight_rom[79] = -14;
        weight_rom[80] = 28;
        weight_rom[81] = 35;
        weight_rom[82] = 3;
        weight_rom[83] = 1;
        weight_rom[84] = 1;
        weight_rom[85] = 2;
        weight_rom[86] = 15;
        weight_rom[87] = -3;
        weight_rom[88] = 0;
        weight_rom[89] = 34;
        weight_rom[90] = -9;
        weight_rom[91] = 0;
        weight_rom[92] = 11;
        weight_rom[93] = 16;
        weight_rom[94] = 41;
        weight_rom[95] = 16;
        weight_rom[96] = 32;
        weight_rom[97] = 48;
        weight_rom[98] = 22;
        weight_rom[99] = 21;
        weight_rom[100] = 30;
        weight_rom[101] = 6;
        weight_rom[102] = 6;
        weight_rom[103] = -12;
        weight_rom[104] = 12;
        weight_rom[105] = 3;
        weight_rom[106] = -10;
        weight_rom[107] = -1;
        weight_rom[108] = -9;
        weight_rom[109] = 45;
        weight_rom[110] = -3;
        weight_rom[111] = -3;
        weight_rom[112] = -1;
        weight_rom[113] = -1;
        weight_rom[114] = 22;
        weight_rom[115] = 0;
        weight_rom[116] = -31;
        weight_rom[117] = 4;
        weight_rom[118] = 47;
        weight_rom[119] = 1;
        weight_rom[120] = 28;
        weight_rom[121] = 34;
        weight_rom[122] = 46;
        weight_rom[123] = 36;
        weight_rom[124] = 39;
        weight_rom[125] = 52;
        weight_rom[126] = 58;
        weight_rom[127] = 45;
        weight_rom[128] = 37;
        weight_rom[129] = 14;
        weight_rom[130] = 30;
        weight_rom[131] = 9;
        weight_rom[132] = 0;
        weight_rom[133] = -26;
        weight_rom[134] = -40;
        weight_rom[135] = -43;
        weight_rom[136] = -19;
        weight_rom[137] = 9;
        weight_rom[138] = 34;
        weight_rom[139] = 1;
        weight_rom[140] = 1;
        weight_rom[141] = 2;
        weight_rom[142] = -2;
        weight_rom[143] = 30;
        weight_rom[144] = 24;
        weight_rom[145] = 10;
        weight_rom[146] = -20;
        weight_rom[147] = 19;
        weight_rom[148] = -10;
        weight_rom[149] = -4;
        weight_rom[150] = 12;
        weight_rom[151] = 17;
        weight_rom[152] = 33;
        weight_rom[153] = 36;
        weight_rom[154] = 24;
        weight_rom[155] = 29;
        weight_rom[156] = 23;
        weight_rom[157] = 6;
        weight_rom[158] = 4;
        weight_rom[159] = 0;
        weight_rom[160] = 4;
        weight_rom[161] = -1;
        weight_rom[162] = -5;
        weight_rom[163] = -28;
        weight_rom[164] = -6;
        weight_rom[165] = 13;
        weight_rom[166] = 17;
        weight_rom[167] = -1;
        weight_rom[168] = -1;
        weight_rom[169] = 3;
        weight_rom[170] = -21;
        weight_rom[171] = 26;
        weight_rom[172] = -43;
        weight_rom[173] = -13;
        weight_rom[174] = -15;
        weight_rom[175] = -10;
        weight_rom[176] = -12;
        weight_rom[177] = 11;
        weight_rom[178] = 12;
        weight_rom[179] = 23;
        weight_rom[180] = 18;
        weight_rom[181] = 35;
        weight_rom[182] = 36;
        weight_rom[183] = 35;
        weight_rom[184] = 35;
        weight_rom[185] = 17;
        weight_rom[186] = 18;
        weight_rom[187] = 7;
        weight_rom[188] = 1;
        weight_rom[189] = -15;
        weight_rom[190] = -20;
        weight_rom[191] = -16;
        weight_rom[192] = 13;
        weight_rom[193] = 40;
        weight_rom[194] = 10;
        weight_rom[195] = 3;
        weight_rom[196] = 0;
        weight_rom[197] = 34;
        weight_rom[198] = -27;
        weight_rom[199] = -22;
        weight_rom[200] = -2;
        weight_rom[201] = -34;
        weight_rom[202] = -20;
        weight_rom[203] = -32;
        weight_rom[204] = 15;
        weight_rom[205] = -9;
        weight_rom[206] = 11;
        weight_rom[207] = 2;
        weight_rom[208] = 21;
        weight_rom[209] = 18;
        weight_rom[210] = 35;
        weight_rom[211] = 34;
        weight_rom[212] = 34;
        weight_rom[213] = 8;
        weight_rom[214] = 16;
        weight_rom[215] = 5;
        weight_rom[216] = 9;
        weight_rom[217] = 0;
        weight_rom[218] = -11;
        weight_rom[219] = -11;
        weight_rom[220] = 7;
        weight_rom[221] = 14;
        weight_rom[222] = 10;
        weight_rom[223] = 19;
        weight_rom[224] = -24;
        weight_rom[225] = -10;
        weight_rom[226] = -34;
        weight_rom[227] = -12;
        weight_rom[228] = 9;
        weight_rom[229] = -12;
        weight_rom[230] = 8;
        weight_rom[231] = 18;
        weight_rom[232] = -9;
        weight_rom[233] = -8;
        weight_rom[234] = 4;
        weight_rom[235] = -8;
        weight_rom[236] = 14;
        weight_rom[237] = 25;
        weight_rom[238] = 33;
        weight_rom[239] = 26;
        weight_rom[240] = 18;
        weight_rom[241] = 11;
        weight_rom[242] = 6;
        weight_rom[243] = 18;
        weight_rom[244] = 7;
        weight_rom[245] = 10;
        weight_rom[246] = 10;
        weight_rom[247] = 7;
        weight_rom[248] = 3;
        weight_rom[249] = 18;
        weight_rom[250] = 71;
        weight_rom[251] = 48;
        weight_rom[252] = -8;
        weight_rom[253] = -9;
        weight_rom[254] = -32;
        weight_rom[255] = 8;
        weight_rom[256] = 13;
        weight_rom[257] = 4;
        weight_rom[258] = 22;
        weight_rom[259] = 10;
        weight_rom[260] = 9;
        weight_rom[261] = 14;
        weight_rom[262] = 5;
        weight_rom[263] = 6;
        weight_rom[264] = 0;
        weight_rom[265] = 1;
        weight_rom[266] = 11;
        weight_rom[267] = 13;
        weight_rom[268] = 1;
        weight_rom[269] = 8;
        weight_rom[270] = 2;
        weight_rom[271] = 13;
        weight_rom[272] = 10;
        weight_rom[273] = 8;
        weight_rom[274] = 25;
        weight_rom[275] = 20;
        weight_rom[276] = 11;
        weight_rom[277] = 55;
        weight_rom[278] = 28;
        weight_rom[279] = -23;
        weight_rom[280] = -18;
        weight_rom[281] = -18;
        weight_rom[282] = -55;
        weight_rom[283] = 9;
        weight_rom[284] = 18;
        weight_rom[285] = 14;
        weight_rom[286] = 31;
        weight_rom[287] = 11;
        weight_rom[288] = 4;
        weight_rom[289] = -2;
        weight_rom[290] = -1;
        weight_rom[291] = 0;
        weight_rom[292] = -5;
        weight_rom[293] = -15;
        weight_rom[294] = -2;
        weight_rom[295] = -11;
        weight_rom[296] = 4;
        weight_rom[297] = 1;
        weight_rom[298] = 8;
        weight_rom[299] = 3;
        weight_rom[300] = 2;
        weight_rom[301] = 17;
        weight_rom[302] = 9;
        weight_rom[303] = 42;
        weight_rom[304] = 30;
        weight_rom[305] = 49;
        weight_rom[306] = 48;
        weight_rom[307] = 31;
        weight_rom[308] = -27;
        weight_rom[309] = -37;
        weight_rom[310] = -35;
        weight_rom[311] = 1;
        weight_rom[312] = 14;
        weight_rom[313] = 19;
        weight_rom[314] = -1;
        weight_rom[315] = -11;
        weight_rom[316] = 6;
        weight_rom[317] = -18;
        weight_rom[318] = -18;
        weight_rom[319] = -13;
        weight_rom[320] = -34;
        weight_rom[321] = 0;
        weight_rom[322] = 15;
        weight_rom[323] = 3;
        weight_rom[324] = -10;
        weight_rom[325] = 0;
        weight_rom[326] = 19;
        weight_rom[327] = 21;
        weight_rom[328] = 10;
        weight_rom[329] = 4;
        weight_rom[330] = 21;
        weight_rom[331] = 15;
        weight_rom[332] = 61;
        weight_rom[333] = 90;
        weight_rom[334] = 70;
        weight_rom[335] = -1;
        weight_rom[336] = -17;
        weight_rom[337] = -21;
        weight_rom[338] = -46;
        weight_rom[339] = 3;
        weight_rom[340] = 27;
        weight_rom[341] = 15;
        weight_rom[342] = -11;
        weight_rom[343] = -24;
        weight_rom[344] = -31;
        weight_rom[345] = -16;
        weight_rom[346] = -18;
        weight_rom[347] = -30;
        weight_rom[348] = -25;
        weight_rom[349] = 8;
        weight_rom[350] = 37;
        weight_rom[351] = 15;
        weight_rom[352] = -1;
        weight_rom[353] = 5;
        weight_rom[354] = 8;
        weight_rom[355] = 23;
        weight_rom[356] = 34;
        weight_rom[357] = 7;
        weight_rom[358] = -6;
        weight_rom[359] = -17;
        weight_rom[360] = 9;
        weight_rom[361] = 64;
        weight_rom[362] = 84;
        weight_rom[363] = 0;
        weight_rom[364] = -2;
        weight_rom[365] = -15;
        weight_rom[366] = -44;
        weight_rom[367] = 32;
        weight_rom[368] = -13;
        weight_rom[369] = -36;
        weight_rom[370] = -42;
        weight_rom[371] = -47;
        weight_rom[372] = -20;
        weight_rom[373] = -19;
        weight_rom[374] = -43;
        weight_rom[375] = -27;
        weight_rom[376] = 10;
        weight_rom[377] = 30;
        weight_rom[378] = 36;
        weight_rom[379] = 22;
        weight_rom[380] = 4;
        weight_rom[381] = -1;
        weight_rom[382] = 2;
        weight_rom[383] = 14;
        weight_rom[384] = 12;
        weight_rom[385] = -6;
        weight_rom[386] = -11;
        weight_rom[387] = -47;
        weight_rom[388] = -41;
        weight_rom[389] = 36;
        weight_rom[390] = 42;
        weight_rom[391] = 2;
        weight_rom[392] = 1;
        weight_rom[393] = -3;
        weight_rom[394] = -11;
        weight_rom[395] = 22;
        weight_rom[396] = -49;
        weight_rom[397] = -42;
        weight_rom[398] = -28;
        weight_rom[399] = -31;
        weight_rom[400] = -18;
        weight_rom[401] = -23;
        weight_rom[402] = -22;
        weight_rom[403] = -20;
        weight_rom[404] = 17;
        weight_rom[405] = 44;
        weight_rom[406] = 36;
        weight_rom[407] = 17;
        weight_rom[408] = 1;
        weight_rom[409] = -4;
        weight_rom[410] = -6;
        weight_rom[411] = -18;
        weight_rom[412] = -12;
        weight_rom[413] = -13;
        weight_rom[414] = -51;
        weight_rom[415] = -60;
        weight_rom[416] = -55;
        weight_rom[417] = -19;
        weight_rom[418] = 51;
        weight_rom[419] = -3;
        weight_rom[420] = -3;
        weight_rom[421] = -9;
        weight_rom[422] = -33;
        weight_rom[423] = 13;
        weight_rom[424] = 6;
        weight_rom[425] = -32;
        weight_rom[426] = -4;
        weight_rom[427] = -11;
        weight_rom[428] = -11;
        weight_rom[429] = -11;
        weight_rom[430] = -17;
        weight_rom[431] = -9;
        weight_rom[432] = 15;
        weight_rom[433] = 49;
        weight_rom[434] = 32;
        weight_rom[435] = 6;
        weight_rom[436] = -4;
        weight_rom[437] = -16;
        weight_rom[438] = -13;
        weight_rom[439] = -21;
        weight_rom[440] = -39;
        weight_rom[441] = -46;
        weight_rom[442] = -47;
        weight_rom[443] = -57;
        weight_rom[444] = -16;
        weight_rom[445] = 10;
        weight_rom[446] = 26;
        weight_rom[447] = 24;
        weight_rom[448] = -2;
        weight_rom[449] = 2;
        weight_rom[450] = 38;
        weight_rom[451] = 67;
        weight_rom[452] = 34;
        weight_rom[453] = 4;
        weight_rom[454] = -5;
        weight_rom[455] = -14;
        weight_rom[456] = -25;
        weight_rom[457] = -4;
        weight_rom[458] = 6;
        weight_rom[459] = 10;
        weight_rom[460] = 33;
        weight_rom[461] = 30;
        weight_rom[462] = 18;
        weight_rom[463] = -8;
        weight_rom[464] = 2;
        weight_rom[465] = -9;
        weight_rom[466] = -17;
        weight_rom[467] = -35;
        weight_rom[468] = -37;
        weight_rom[469] = -32;
        weight_rom[470] = -15;
        weight_rom[471] = 0;
        weight_rom[472] = 20;
        weight_rom[473] = 47;
        weight_rom[474] = 56;
        weight_rom[475] = 43;
        weight_rom[476] = 2;
        weight_rom[477] = 0;
        weight_rom[478] = 7;
        weight_rom[479] = 67;
        weight_rom[480] = 32;
        weight_rom[481] = 5;
        weight_rom[482] = 13;
        weight_rom[483] = 2;
        weight_rom[484] = 1;
        weight_rom[485] = 5;
        weight_rom[486] = 14;
        weight_rom[487] = 27;
        weight_rom[488] = 34;
        weight_rom[489] = 14;
        weight_rom[490] = -3;
        weight_rom[491] = -9;
        weight_rom[492] = -2;
        weight_rom[493] = -14;
        weight_rom[494] = -25;
        weight_rom[495] = -10;
        weight_rom[496] = -24;
        weight_rom[497] = -16;
        weight_rom[498] = -14;
        weight_rom[499] = 16;
        weight_rom[500] = 20;
        weight_rom[501] = 9;
        weight_rom[502] = 60;
        weight_rom[503] = -1;
        weight_rom[504] = 1;
        weight_rom[505] = -1;
        weight_rom[506] = 46;
        weight_rom[507] = 27;
        weight_rom[508] = 1;
        weight_rom[509] = 11;
        weight_rom[510] = 17;
        weight_rom[511] = -11;
        weight_rom[512] = -4;
        weight_rom[513] = 3;
        weight_rom[514] = 17;
        weight_rom[515] = 21;
        weight_rom[516] = 14;
        weight_rom[517] = 6;
        weight_rom[518] = -3;
        weight_rom[519] = -2;
        weight_rom[520] = -1;
        weight_rom[521] = -3;
        weight_rom[522] = 3;
        weight_rom[523] = 2;
        weight_rom[524] = 5;
        weight_rom[525] = -7;
        weight_rom[526] = 17;
        weight_rom[527] = 32;
        weight_rom[528] = 53;
        weight_rom[529] = 39;
        weight_rom[530] = 29;
        weight_rom[531] = 36;
        weight_rom[532] = -1;
        weight_rom[533] = 2;
        weight_rom[534] = -22;
        weight_rom[535] = -14;
        weight_rom[536] = 6;
        weight_rom[537] = 12;
        weight_rom[538] = 4;
        weight_rom[539] = 22;
        weight_rom[540] = 19;
        weight_rom[541] = 26;
        weight_rom[542] = 13;
        weight_rom[543] = -8;
        weight_rom[544] = -7;
        weight_rom[545] = -2;
        weight_rom[546] = -3;
        weight_rom[547] = -1;
        weight_rom[548] = 1;
        weight_rom[549] = 8;
        weight_rom[550] = 12;
        weight_rom[551] = 5;
        weight_rom[552] = 3;
        weight_rom[553] = 6;
        weight_rom[554] = 36;
        weight_rom[555] = 53;
        weight_rom[556] = 31;
        weight_rom[557] = 31;
        weight_rom[558] = 36;
        weight_rom[559] = 16;
        weight_rom[560] = 0;
        weight_rom[561] = -23;
        weight_rom[562] = -23;
        weight_rom[563] = 6;
        weight_rom[564] = 26;
        weight_rom[565] = 20;
        weight_rom[566] = 36;
        weight_rom[567] = 47;
        weight_rom[568] = 35;
        weight_rom[569] = 20;
        weight_rom[570] = 18;
        weight_rom[571] = -5;
        weight_rom[572] = -9;
        weight_rom[573] = -18;
        weight_rom[574] = -20;
        weight_rom[575] = -15;
        weight_rom[576] = -1;
        weight_rom[577] = 4;
        weight_rom[578] = 14;
        weight_rom[579] = 18;
        weight_rom[580] = 24;
        weight_rom[581] = 43;
        weight_rom[582] = 41;
        weight_rom[583] = 48;
        weight_rom[584] = 24;
        weight_rom[585] = 31;
        weight_rom[586] = 10;
        weight_rom[587] = 2;
        weight_rom[588] = -2;
        weight_rom[589] = 12;
        weight_rom[590] = 35;
        weight_rom[591] = 60;
        weight_rom[592] = 47;
        weight_rom[593] = 29;
        weight_rom[594] = 56;
        weight_rom[595] = 42;
        weight_rom[596] = 31;
        weight_rom[597] = 14;
        weight_rom[598] = -2;
        weight_rom[599] = -5;
        weight_rom[600] = -22;
        weight_rom[601] = -6;
        weight_rom[602] = -7;
        weight_rom[603] = -12;
        weight_rom[604] = -3;
        weight_rom[605] = 3;
        weight_rom[606] = 16;
        weight_rom[607] = 34;
        weight_rom[608] = 17;
        weight_rom[609] = 37;
        weight_rom[610] = 37;
        weight_rom[611] = 20;
        weight_rom[612] = 47;
        weight_rom[613] = 41;
        weight_rom[614] = -24;
        weight_rom[615] = 2;
        weight_rom[616] = 0;
        weight_rom[617] = 1;
        weight_rom[618] = 24;
        weight_rom[619] = 48;
        weight_rom[620] = 43;
        weight_rom[621] = 53;
        weight_rom[622] = 44;
        weight_rom[623] = 34;
        weight_rom[624] = 11;
        weight_rom[625] = 1;
        weight_rom[626] = 5;
        weight_rom[627] = 8;
        weight_rom[628] = -4;
        weight_rom[629] = -7;
        weight_rom[630] = 18;
        weight_rom[631] = 9;
        weight_rom[632] = 3;
        weight_rom[633] = 23;
        weight_rom[634] = 22;
        weight_rom[635] = 18;
        weight_rom[636] = 25;
        weight_rom[637] = 13;
        weight_rom[638] = 10;
        weight_rom[639] = 8;
        weight_rom[640] = 50;
        weight_rom[641] = 35;
        weight_rom[642] = 11;
        weight_rom[643] = -1;
        weight_rom[644] = 2;
        weight_rom[645] = 2;
        weight_rom[646] = 27;
        weight_rom[647] = 19;
        weight_rom[648] = 28;
        weight_rom[649] = 6;
        weight_rom[650] = 6;
        weight_rom[651] = -5;
        weight_rom[652] = 26;
        weight_rom[653] = 21;
        weight_rom[654] = 18;
        weight_rom[655] = 27;
        weight_rom[656] = 37;
        weight_rom[657] = 39;
        weight_rom[658] = 16;
        weight_rom[659] = 19;
        weight_rom[660] = 24;
        weight_rom[661] = 9;
        weight_rom[662] = 5;
        weight_rom[663] = 25;
        weight_rom[664] = 24;
        weight_rom[665] = -12;
        weight_rom[666] = 28;
        weight_rom[667] = 27;
        weight_rom[668] = 10;
        weight_rom[669] = -8;
        weight_rom[670] = 28;
        weight_rom[671] = 3;
        weight_rom[672] = 2;
        weight_rom[673] = 0;
        weight_rom[674] = 20;
        weight_rom[675] = -34;
        weight_rom[676] = -1;
        weight_rom[677] = -37;
        weight_rom[678] = -26;
        weight_rom[679] = -9;
        weight_rom[680] = -9;
        weight_rom[681] = 16;
        weight_rom[682] = 7;
        weight_rom[683] = 22;
        weight_rom[684] = 32;
        weight_rom[685] = 22;
        weight_rom[686] = 26;
        weight_rom[687] = 24;
        weight_rom[688] = 12;
        weight_rom[689] = 12;
        weight_rom[690] = 40;
        weight_rom[691] = 33;
        weight_rom[692] = 28;
        weight_rom[693] = 47;
        weight_rom[694] = 20;
        weight_rom[695] = 31;
        weight_rom[696] = 25;
        weight_rom[697] = 30;
        weight_rom[698] = 1;
        weight_rom[699] = -1;
        weight_rom[700] = -3;
        weight_rom[701] = -2;
        weight_rom[702] = -2;
        weight_rom[703] = -24;
        weight_rom[704] = -30;
        weight_rom[705] = -31;
        weight_rom[706] = -2;
        weight_rom[707] = 5;
        weight_rom[708] = 18;
        weight_rom[709] = 9;
        weight_rom[710] = 12;
        weight_rom[711] = 10;
        weight_rom[712] = 25;
        weight_rom[713] = 11;
        weight_rom[714] = 29;
        weight_rom[715] = 13;
        weight_rom[716] = 38;
        weight_rom[717] = 41;
        weight_rom[718] = 38;
        weight_rom[719] = 43;
        weight_rom[720] = 58;
        weight_rom[721] = 43;
        weight_rom[722] = 3;
        weight_rom[723] = 25;
        weight_rom[724] = 32;
        weight_rom[725] = -3;
        weight_rom[726] = 2;
        weight_rom[727] = 1;
        weight_rom[728] = 0;
        weight_rom[729] = -1;
        weight_rom[730] = 2;
        weight_rom[731] = 1;
        weight_rom[732] = -3;
        weight_rom[733] = -12;
        weight_rom[734] = 9;
        weight_rom[735] = 15;
        weight_rom[736] = 19;
        weight_rom[737] = 53;
        weight_rom[738] = 35;
        weight_rom[739] = 37;
        weight_rom[740] = 43;
        weight_rom[741] = 48;
        weight_rom[742] = 67;
        weight_rom[743] = 36;
        weight_rom[744] = 48;
        weight_rom[745] = 59;
        weight_rom[746] = 52;
        weight_rom[747] = 33;
        weight_rom[748] = 46;
        weight_rom[749] = 40;
        weight_rom[750] = 19;
        weight_rom[751] = 38;
        weight_rom[752] = -1;
        weight_rom[753] = 2;
        weight_rom[754] = -1;
        weight_rom[755] = -1;
        weight_rom[756] = -3;
        weight_rom[757] = 3;
        weight_rom[758] = -1;
        weight_rom[759] = -1;
        weight_rom[760] = -1;
        weight_rom[761] = -21;
        weight_rom[762] = -40;
        weight_rom[763] = -26;
        weight_rom[764] = -38;
        weight_rom[765] = -1;
        weight_rom[766] = -10;
        weight_rom[767] = 24;
        weight_rom[768] = 4;
        weight_rom[769] = -50;
        weight_rom[770] = 35;
        weight_rom[771] = -20;
        weight_rom[772] = -16;
        weight_rom[773] = -67;
        weight_rom[774] = -40;
        weight_rom[775] = -17;
        weight_rom[776] = -7;
        weight_rom[777] = 17;
        weight_rom[778] = 20;
        weight_rom[779] = -1;
        weight_rom[780] = -2;
        weight_rom[781] = 2;
        weight_rom[782] = 3;
        weight_rom[783] = 1;
        weight_rom[784] = -1;
        weight_rom[785] = 2;
        weight_rom[786] = 0;
        weight_rom[787] = 0;
        weight_rom[788] = 0;
        weight_rom[789] = 0;
        weight_rom[790] = 1;
        weight_rom[791] = 1;
        weight_rom[792] = 1;
        weight_rom[793] = -3;
        weight_rom[794] = 2;
        weight_rom[795] = -1;
        weight_rom[796] = -2;
        weight_rom[797] = 12;
        weight_rom[798] = 26;
        weight_rom[799] = -1;
        weight_rom[800] = 2;
        weight_rom[801] = 2;
        weight_rom[802] = -1;
        weight_rom[803] = 3;
        weight_rom[804] = -1;
        weight_rom[805] = 3;
        weight_rom[806] = 1;
        weight_rom[807] = -1;
        weight_rom[808] = 0;
        weight_rom[809] = -1;
        weight_rom[810] = 0;
        weight_rom[811] = 0;
        weight_rom[812] = -3;
        weight_rom[813] = -1;
        weight_rom[814] = 2;
        weight_rom[815] = 1;
        weight_rom[816] = 2;
        weight_rom[817] = 0;
        weight_rom[818] = -26;
        weight_rom[819] = -33;
        weight_rom[820] = -28;
        weight_rom[821] = -52;
        weight_rom[822] = -53;
        weight_rom[823] = -50;
        weight_rom[824] = -66;
        weight_rom[825] = -56;
        weight_rom[826] = -3;
        weight_rom[827] = -5;
        weight_rom[828] = 43;
        weight_rom[829] = -18;
        weight_rom[830] = -57;
        weight_rom[831] = -39;
        weight_rom[832] = -37;
        weight_rom[833] = -33;
        weight_rom[834] = -37;
        weight_rom[835] = -22;
        weight_rom[836] = -3;
        weight_rom[837] = -2;
        weight_rom[838] = -1;
        weight_rom[839] = 2;
        weight_rom[840] = 1;
        weight_rom[841] = 1;
        weight_rom[842] = 1;
        weight_rom[843] = 0;
        weight_rom[844] = -19;
        weight_rom[845] = -2;
        weight_rom[846] = -40;
        weight_rom[847] = -50;
        weight_rom[848] = -26;
        weight_rom[849] = 10;
        weight_rom[850] = -39;
        weight_rom[851] = -13;
        weight_rom[852] = -27;
        weight_rom[853] = -7;
        weight_rom[854] = -14;
        weight_rom[855] = -18;
        weight_rom[856] = -3;
        weight_rom[857] = -20;
        weight_rom[858] = -32;
        weight_rom[859] = -33;
        weight_rom[860] = -20;
        weight_rom[861] = -15;
        weight_rom[862] = -31;
        weight_rom[863] = -10;
        weight_rom[864] = -18;
        weight_rom[865] = -20;
        weight_rom[866] = 2;
        weight_rom[867] = 1;
        weight_rom[868] = -3;
        weight_rom[869] = -2;
        weight_rom[870] = -19;
        weight_rom[871] = 0;
        weight_rom[872] = 2;
        weight_rom[873] = 7;
        weight_rom[874] = -37;
        weight_rom[875] = -25;
        weight_rom[876] = -20;
        weight_rom[877] = -14;
        weight_rom[878] = -8;
        weight_rom[879] = 6;
        weight_rom[880] = -3;
        weight_rom[881] = -15;
        weight_rom[882] = -7;
        weight_rom[883] = -29;
        weight_rom[884] = -13;
        weight_rom[885] = -2;
        weight_rom[886] = -8;
        weight_rom[887] = -13;
        weight_rom[888] = -20;
        weight_rom[889] = -41;
        weight_rom[890] = -37;
        weight_rom[891] = -49;
        weight_rom[892] = -44;
        weight_rom[893] = -21;
        weight_rom[894] = -1;
        weight_rom[895] = -2;
        weight_rom[896] = 0;
        weight_rom[897] = 2;
        weight_rom[898] = 9;
        weight_rom[899] = 1;
        weight_rom[900] = -31;
        weight_rom[901] = -3;
        weight_rom[902] = 22;
        weight_rom[903] = 3;
        weight_rom[904] = 17;
        weight_rom[905] = 10;
        weight_rom[906] = 13;
        weight_rom[907] = 13;
        weight_rom[908] = 18;
        weight_rom[909] = 15;
        weight_rom[910] = 10;
        weight_rom[911] = 4;
        weight_rom[912] = -4;
        weight_rom[913] = -4;
        weight_rom[914] = -1;
        weight_rom[915] = -21;
        weight_rom[916] = 4;
        weight_rom[917] = -33;
        weight_rom[918] = -26;
        weight_rom[919] = -48;
        weight_rom[920] = -62;
        weight_rom[921] = -11;
        weight_rom[922] = 2;
        weight_rom[923] = 3;
        weight_rom[924] = 1;
        weight_rom[925] = -2;
        weight_rom[926] = 1;
        weight_rom[927] = 26;
        weight_rom[928] = 46;
        weight_rom[929] = 35;
        weight_rom[930] = 17;
        weight_rom[931] = 20;
        weight_rom[932] = 21;
        weight_rom[933] = 27;
        weight_rom[934] = 8;
        weight_rom[935] = 21;
        weight_rom[936] = 19;
        weight_rom[937] = 20;
        weight_rom[938] = 14;
        weight_rom[939] = 10;
        weight_rom[940] = 17;
        weight_rom[941] = 6;
        weight_rom[942] = 1;
        weight_rom[943] = -11;
        weight_rom[944] = -21;
        weight_rom[945] = -25;
        weight_rom[946] = -18;
        weight_rom[947] = -25;
        weight_rom[948] = -15;
        weight_rom[949] = -3;
        weight_rom[950] = -18;
        weight_rom[951] = -1;
        weight_rom[952] = 3;
        weight_rom[953] = 2;
        weight_rom[954] = -9;
        weight_rom[955] = 59;
        weight_rom[956] = 30;
        weight_rom[957] = 14;
        weight_rom[958] = 40;
        weight_rom[959] = 20;
        weight_rom[960] = 21;
        weight_rom[961] = 24;
        weight_rom[962] = 28;
        weight_rom[963] = 16;
        weight_rom[964] = 13;
        weight_rom[965] = 22;
        weight_rom[966] = 28;
        weight_rom[967] = 22;
        weight_rom[968] = 30;
        weight_rom[969] = 15;
        weight_rom[970] = 10;
        weight_rom[971] = -6;
        weight_rom[972] = -8;
        weight_rom[973] = -8;
        weight_rom[974] = -13;
        weight_rom[975] = -48;
        weight_rom[976] = -65;
        weight_rom[977] = -36;
        weight_rom[978] = -15;
        weight_rom[979] = 17;
        weight_rom[980] = -2;
        weight_rom[981] = -6;
        weight_rom[982] = 63;
        weight_rom[983] = 60;
        weight_rom[984] = 34;
        weight_rom[985] = 18;
        weight_rom[986] = 32;
        weight_rom[987] = 19;
        weight_rom[988] = 8;
        weight_rom[989] = 12;
        weight_rom[990] = 15;
        weight_rom[991] = 8;
        weight_rom[992] = 8;
        weight_rom[993] = 17;
        weight_rom[994] = 20;
        weight_rom[995] = 20;
        weight_rom[996] = 23;
        weight_rom[997] = 13;
        weight_rom[998] = 8;
        weight_rom[999] = 7;
        weight_rom[1000] = 1;
        weight_rom[1001] = -5;
        weight_rom[1002] = -4;
        weight_rom[1003] = -29;
        weight_rom[1004] = -45;
        weight_rom[1005] = -43;
        weight_rom[1006] = -10;
        weight_rom[1007] = -2;
        weight_rom[1008] = 17;
        weight_rom[1009] = 27;
        weight_rom[1010] = 16;
        weight_rom[1011] = 43;
        weight_rom[1012] = 43;
        weight_rom[1013] = 20;
        weight_rom[1014] = 21;
        weight_rom[1015] = 25;
        weight_rom[1016] = 23;
        weight_rom[1017] = 9;
        weight_rom[1018] = 17;
        weight_rom[1019] = 12;
        weight_rom[1020] = 13;
        weight_rom[1021] = 10;
        weight_rom[1022] = 25;
        weight_rom[1023] = 29;
        weight_rom[1024] = 23;
        weight_rom[1025] = 21;
        weight_rom[1026] = 18;
        weight_rom[1027] = 16;
        weight_rom[1028] = 12;
        weight_rom[1029] = 1;
        weight_rom[1030] = 12;
        weight_rom[1031] = -18;
        weight_rom[1032] = -70;
        weight_rom[1033] = -37;
        weight_rom[1034] = -40;
        weight_rom[1035] = -17;
        weight_rom[1036] = 21;
        weight_rom[1037] = 37;
        weight_rom[1038] = 29;
        weight_rom[1039] = 51;
        weight_rom[1040] = 57;
        weight_rom[1041] = 38;
        weight_rom[1042] = 14;
        weight_rom[1043] = 7;
        weight_rom[1044] = -3;
        weight_rom[1045] = -2;
        weight_rom[1046] = 2;
        weight_rom[1047] = -4;
        weight_rom[1048] = -1;
        weight_rom[1049] = 6;
        weight_rom[1050] = 20;
        weight_rom[1051] = 22;
        weight_rom[1052] = 28;
        weight_rom[1053] = 28;
        weight_rom[1054] = 23;
        weight_rom[1055] = 22;
        weight_rom[1056] = 16;
        weight_rom[1057] = -3;
        weight_rom[1058] = 7;
        weight_rom[1059] = -10;
        weight_rom[1060] = -49;
        weight_rom[1061] = -65;
        weight_rom[1062] = -25;
        weight_rom[1063] = 17;
        weight_rom[1064] = 24;
        weight_rom[1065] = 42;
        weight_rom[1066] = 54;
        weight_rom[1067] = 50;
        weight_rom[1068] = 7;
        weight_rom[1069] = 24;
        weight_rom[1070] = 16;
        weight_rom[1071] = -10;
        weight_rom[1072] = -13;
        weight_rom[1073] = -14;
        weight_rom[1074] = -15;
        weight_rom[1075] = -24;
        weight_rom[1076] = -27;
        weight_rom[1077] = -16;
        weight_rom[1078] = 1;
        weight_rom[1079] = 13;
        weight_rom[1080] = 30;
        weight_rom[1081] = 30;
        weight_rom[1082] = 33;
        weight_rom[1083] = 40;
        weight_rom[1084] = 29;
        weight_rom[1085] = 26;
        weight_rom[1086] = 34;
        weight_rom[1087] = -1;
        weight_rom[1088] = -58;
        weight_rom[1089] = -85;
        weight_rom[1090] = -39;
        weight_rom[1091] = -13;
        weight_rom[1092] = 19;
        weight_rom[1093] = 61;
        weight_rom[1094] = 74;
        weight_rom[1095] = 50;
        weight_rom[1096] = 15;
        weight_rom[1097] = 4;
        weight_rom[1098] = -17;
        weight_rom[1099] = -5;
        weight_rom[1100] = -27;
        weight_rom[1101] = -20;
        weight_rom[1102] = -19;
        weight_rom[1103] = -19;
        weight_rom[1104] = -27;
        weight_rom[1105] = -46;
        weight_rom[1106] = -22;
        weight_rom[1107] = 3;
        weight_rom[1108] = 13;
        weight_rom[1109] = 18;
        weight_rom[1110] = 31;
        weight_rom[1111] = 31;
        weight_rom[1112] = 39;
        weight_rom[1113] = 31;
        weight_rom[1114] = 43;
        weight_rom[1115] = 10;
        weight_rom[1116] = -44;
        weight_rom[1117] = -60;
        weight_rom[1118] = -72;
        weight_rom[1119] = -24;
        weight_rom[1120] = 10;
        weight_rom[1121] = 34;
        weight_rom[1122] = 71;
        weight_rom[1123] = 48;
        weight_rom[1124] = 2;
        weight_rom[1125] = -15;
        weight_rom[1126] = -32;
        weight_rom[1127] = -23;
        weight_rom[1128] = -13;
        weight_rom[1129] = -19;
        weight_rom[1130] = -27;
        weight_rom[1131] = -21;
        weight_rom[1132] = -28;
        weight_rom[1133] = -59;
        weight_rom[1134] = -26;
        weight_rom[1135] = -8;
        weight_rom[1136] = 12;
        weight_rom[1137] = 9;
        weight_rom[1138] = 21;
        weight_rom[1139] = 21;
        weight_rom[1140] = 17;
        weight_rom[1141] = 12;
        weight_rom[1142] = 13;
        weight_rom[1143] = -3;
        weight_rom[1144] = -9;
        weight_rom[1145] = -5;
        weight_rom[1146] = 26;
        weight_rom[1147] = -26;
        weight_rom[1148] = 2;
        weight_rom[1149] = 9;
        weight_rom[1150] = 72;
        weight_rom[1151] = 3;
        weight_rom[1152] = -2;
        weight_rom[1153] = -30;
        weight_rom[1154] = -23;
        weight_rom[1155] = -21;
        weight_rom[1156] = -14;
        weight_rom[1157] = -1;
        weight_rom[1158] = 0;
        weight_rom[1159] = -9;
        weight_rom[1160] = -36;
        weight_rom[1161] = -32;
        weight_rom[1162] = -13;
        weight_rom[1163] = -6;
        weight_rom[1164] = 12;
        weight_rom[1165] = 10;
        weight_rom[1166] = 8;
        weight_rom[1167] = 3;
        weight_rom[1168] = 8;
        weight_rom[1169] = -3;
        weight_rom[1170] = -11;
        weight_rom[1171] = 2;
        weight_rom[1172] = 1;
        weight_rom[1173] = 40;
        weight_rom[1174] = 47;
        weight_rom[1175] = 40;
        weight_rom[1176] = -1;
        weight_rom[1177] = 26;
        weight_rom[1178] = 25;
        weight_rom[1179] = -5;
        weight_rom[1180] = -27;
        weight_rom[1181] = -12;
        weight_rom[1182] = -14;
        weight_rom[1183] = 5;
        weight_rom[1184] = -4;
        weight_rom[1185] = -6;
        weight_rom[1186] = -7;
        weight_rom[1187] = -9;
        weight_rom[1188] = -16;
        weight_rom[1189] = -25;
        weight_rom[1190] = -6;
        weight_rom[1191] = -5;
        weight_rom[1192] = 0;
        weight_rom[1193] = 14;
        weight_rom[1194] = 26;
        weight_rom[1195] = 27;
        weight_rom[1196] = 18;
        weight_rom[1197] = 0;
        weight_rom[1198] = 2;
        weight_rom[1199] = 22;
        weight_rom[1200] = -16;
        weight_rom[1201] = 30;
        weight_rom[1202] = 68;
        weight_rom[1203] = -2;
        weight_rom[1204] = 1;
        weight_rom[1205] = -25;
        weight_rom[1206] = 4;
        weight_rom[1207] = 5;
        weight_rom[1208] = 14;
        weight_rom[1209] = 6;
        weight_rom[1210] = 13;
        weight_rom[1211] = 8;
        weight_rom[1212] = 3;
        weight_rom[1213] = 1;
        weight_rom[1214] = 1;
        weight_rom[1215] = -7;
        weight_rom[1216] = -18;
        weight_rom[1217] = -14;
        weight_rom[1218] = -6;
        weight_rom[1219] = 5;
        weight_rom[1220] = 6;
        weight_rom[1221] = 26;
        weight_rom[1222] = 16;
        weight_rom[1223] = 14;
        weight_rom[1224] = 3;
        weight_rom[1225] = 16;
        weight_rom[1226] = 15;
        weight_rom[1227] = 0;
        weight_rom[1228] = 31;
        weight_rom[1229] = 16;
        weight_rom[1230] = 68;
        weight_rom[1231] = 23;
        weight_rom[1232] = -3;
        weight_rom[1233] = 2;
        weight_rom[1234] = 0;
        weight_rom[1235] = 15;
        weight_rom[1236] = 26;
        weight_rom[1237] = 14;
        weight_rom[1238] = 20;
        weight_rom[1239] = 26;
        weight_rom[1240] = 8;
        weight_rom[1241] = 15;
        weight_rom[1242] = 10;
        weight_rom[1243] = -5;
        weight_rom[1244] = 4;
        weight_rom[1245] = -2;
        weight_rom[1246] = -7;
        weight_rom[1247] = 7;
        weight_rom[1248] = 15;
        weight_rom[1249] = 30;
        weight_rom[1250] = 22;
        weight_rom[1251] = 12;
        weight_rom[1252] = 12;
        weight_rom[1253] = 17;
        weight_rom[1254] = 12;
        weight_rom[1255] = 4;
        weight_rom[1256] = 2;
        weight_rom[1257] = 59;
        weight_rom[1258] = 103;
        weight_rom[1259] = 53;
        weight_rom[1260] = 2;
        weight_rom[1261] = -1;
        weight_rom[1262] = 5;
        weight_rom[1263] = 19;
        weight_rom[1264] = 16;
        weight_rom[1265] = 5;
        weight_rom[1266] = 5;
        weight_rom[1267] = 8;
        weight_rom[1268] = 13;
        weight_rom[1269] = 16;
        weight_rom[1270] = 6;
        weight_rom[1271] = 13;
        weight_rom[1272] = 13;
        weight_rom[1273] = 8;
        weight_rom[1274] = -3;
        weight_rom[1275] = 9;
        weight_rom[1276] = 12;
        weight_rom[1277] = 15;
        weight_rom[1278] = 13;
        weight_rom[1279] = 10;
        weight_rom[1280] = 4;
        weight_rom[1281] = 4;
        weight_rom[1282] = 13;
        weight_rom[1283] = 11;
        weight_rom[1284] = 12;
        weight_rom[1285] = 85;
        weight_rom[1286] = 92;
        weight_rom[1287] = -2;
        weight_rom[1288] = -2;
        weight_rom[1289] = -1;
        weight_rom[1290] = 16;
        weight_rom[1291] = -17;
        weight_rom[1292] = 16;
        weight_rom[1293] = 25;
        weight_rom[1294] = -6;
        weight_rom[1295] = 16;
        weight_rom[1296] = 7;
        weight_rom[1297] = 7;
        weight_rom[1298] = 7;
        weight_rom[1299] = 5;
        weight_rom[1300] = -4;
        weight_rom[1301] = 7;
        weight_rom[1302] = 1;
        weight_rom[1303] = 5;
        weight_rom[1304] = 16;
        weight_rom[1305] = 21;
        weight_rom[1306] = 19;
        weight_rom[1307] = 14;
        weight_rom[1308] = -1;
        weight_rom[1309] = 0;
        weight_rom[1310] = -3;
        weight_rom[1311] = -9;
        weight_rom[1312] = 13;
        weight_rom[1313] = 52;
        weight_rom[1314] = 22;
        weight_rom[1315] = 34;
        weight_rom[1316] = 3;
        weight_rom[1317] = -1;
        weight_rom[1318] = -19;
        weight_rom[1319] = 14;
        weight_rom[1320] = 1;
        weight_rom[1321] = 6;
        weight_rom[1322] = 3;
        weight_rom[1323] = 10;
        weight_rom[1324] = 8;
        weight_rom[1325] = 7;
        weight_rom[1326] = -6;
        weight_rom[1327] = -12;
        weight_rom[1328] = -7;
        weight_rom[1329] = -4;
        weight_rom[1330] = 0;
        weight_rom[1331] = -7;
        weight_rom[1332] = -3;
        weight_rom[1333] = 7;
        weight_rom[1334] = -12;
        weight_rom[1335] = -4;
        weight_rom[1336] = -4;
        weight_rom[1337] = 0;
        weight_rom[1338] = 5;
        weight_rom[1339] = 0;
        weight_rom[1340] = 1;
        weight_rom[1341] = 57;
        weight_rom[1342] = 61;
        weight_rom[1343] = 19;
        weight_rom[1344] = 1;
        weight_rom[1345] = -5;
        weight_rom[1346] = -4;
        weight_rom[1347] = -4;
        weight_rom[1348] = 16;
        weight_rom[1349] = 10;
        weight_rom[1350] = 14;
        weight_rom[1351] = 13;
        weight_rom[1352] = 8;
        weight_rom[1353] = -2;
        weight_rom[1354] = -8;
        weight_rom[1355] = -5;
        weight_rom[1356] = -5;
        weight_rom[1357] = -11;
        weight_rom[1358] = 2;
        weight_rom[1359] = -5;
        weight_rom[1360] = -6;
        weight_rom[1361] = -9;
        weight_rom[1362] = -12;
        weight_rom[1363] = 0;
        weight_rom[1364] = 0;
        weight_rom[1365] = -4;
        weight_rom[1366] = -14;
        weight_rom[1367] = -16;
        weight_rom[1368] = 42;
        weight_rom[1369] = 31;
        weight_rom[1370] = 21;
        weight_rom[1371] = 1;
        weight_rom[1372] = -1;
        weight_rom[1373] = 4;
        weight_rom[1374] = 23;
        weight_rom[1375] = 11;
        weight_rom[1376] = -4;
        weight_rom[1377] = -5;
        weight_rom[1378] = 11;
        weight_rom[1379] = -2;
        weight_rom[1380] = -6;
        weight_rom[1381] = -4;
        weight_rom[1382] = -3;
        weight_rom[1383] = -4;
        weight_rom[1384] = -9;
        weight_rom[1385] = -13;
        weight_rom[1386] = -10;
        weight_rom[1387] = -12;
        weight_rom[1388] = 0;
        weight_rom[1389] = -6;
        weight_rom[1390] = 0;
        weight_rom[1391] = 2;
        weight_rom[1392] = -7;
        weight_rom[1393] = -2;
        weight_rom[1394] = -8;
        weight_rom[1395] = 15;
        weight_rom[1396] = 22;
        weight_rom[1397] = 25;
        weight_rom[1398] = 12;
        weight_rom[1399] = 1;
        weight_rom[1400] = -2;
        weight_rom[1401] = -1;
        weight_rom[1402] = -6;
        weight_rom[1403] = 13;
        weight_rom[1404] = -16;
        weight_rom[1405] = 1;
        weight_rom[1406] = 13;
        weight_rom[1407] = 7;
        weight_rom[1408] = 12;
        weight_rom[1409] = 16;
        weight_rom[1410] = 2;
        weight_rom[1411] = 1;
        weight_rom[1412] = 3;
        weight_rom[1413] = -5;
        weight_rom[1414] = 0;
        weight_rom[1415] = -3;
        weight_rom[1416] = -9;
        weight_rom[1417] = -6;
        weight_rom[1418] = -11;
        weight_rom[1419] = 8;
        weight_rom[1420] = -5;
        weight_rom[1421] = -9;
        weight_rom[1422] = 17;
        weight_rom[1423] = 4;
        weight_rom[1424] = 14;
        weight_rom[1425] = -3;
        weight_rom[1426] = 16;
        weight_rom[1427] = 0;
        weight_rom[1428] = -3;
        weight_rom[1429] = -2;
        weight_rom[1430] = -22;
        weight_rom[1431] = -55;
        weight_rom[1432] = -2;
        weight_rom[1433] = -10;
        weight_rom[1434] = 4;
        weight_rom[1435] = 22;
        weight_rom[1436] = -1;
        weight_rom[1437] = 2;
        weight_rom[1438] = 10;
        weight_rom[1439] = 11;
        weight_rom[1440] = 15;
        weight_rom[1441] = 14;
        weight_rom[1442] = 5;
        weight_rom[1443] = 4;
        weight_rom[1444] = -21;
        weight_rom[1445] = -17;
        weight_rom[1446] = -6;
        weight_rom[1447] = -18;
        weight_rom[1448] = -18;
        weight_rom[1449] = 3;
        weight_rom[1450] = 19;
        weight_rom[1451] = -5;
        weight_rom[1452] = 14;
        weight_rom[1453] = -3;
        weight_rom[1454] = 17;
        weight_rom[1455] = 2;
        weight_rom[1456] = -1;
        weight_rom[1457] = -1;
        weight_rom[1458] = -18;
        weight_rom[1459] = -24;
        weight_rom[1460] = -12;
        weight_rom[1461] = 36;
        weight_rom[1462] = 11;
        weight_rom[1463] = 6;
        weight_rom[1464] = 11;
        weight_rom[1465] = -3;
        weight_rom[1466] = 9;
        weight_rom[1467] = 3;
        weight_rom[1468] = 6;
        weight_rom[1469] = 13;
        weight_rom[1470] = 3;
        weight_rom[1471] = -4;
        weight_rom[1472] = -1;
        weight_rom[1473] = 1;
        weight_rom[1474] = -20;
        weight_rom[1475] = -19;
        weight_rom[1476] = -5;
        weight_rom[1477] = -6;
        weight_rom[1478] = 4;
        weight_rom[1479] = -50;
        weight_rom[1480] = 14;
        weight_rom[1481] = 35;
        weight_rom[1482] = 0;
        weight_rom[1483] = 2;
        weight_rom[1484] = 2;
        weight_rom[1485] = 1;
        weight_rom[1486] = -1;
        weight_rom[1487] = -22;
        weight_rom[1488] = 4;
        weight_rom[1489] = 8;
        weight_rom[1490] = -14;
        weight_rom[1491] = -1;
        weight_rom[1492] = 13;
        weight_rom[1493] = 9;
        weight_rom[1494] = -5;
        weight_rom[1495] = 14;
        weight_rom[1496] = 10;
        weight_rom[1497] = 14;
        weight_rom[1498] = 22;
        weight_rom[1499] = 26;
        weight_rom[1500] = 6;
        weight_rom[1501] = -14;
        weight_rom[1502] = -4;
        weight_rom[1503] = -21;
        weight_rom[1504] = -39;
        weight_rom[1505] = -36;
        weight_rom[1506] = -42;
        weight_rom[1507] = -66;
        weight_rom[1508] = -39;
        weight_rom[1509] = 0;
        weight_rom[1510] = -1;
        weight_rom[1511] = -2;
        weight_rom[1512] = -1;
        weight_rom[1513] = -1;
        weight_rom[1514] = 0;
        weight_rom[1515] = 3;
        weight_rom[1516] = -11;
        weight_rom[1517] = -16;
        weight_rom[1518] = -3;
        weight_rom[1519] = 24;
        weight_rom[1520] = 26;
        weight_rom[1521] = 18;
        weight_rom[1522] = 13;
        weight_rom[1523] = 19;
        weight_rom[1524] = -1;
        weight_rom[1525] = 12;
        weight_rom[1526] = 26;
        weight_rom[1527] = 18;
        weight_rom[1528] = 26;
        weight_rom[1529] = 27;
        weight_rom[1530] = 4;
        weight_rom[1531] = 7;
        weight_rom[1532] = -24;
        weight_rom[1533] = -23;
        weight_rom[1534] = 28;
        weight_rom[1535] = -18;
        weight_rom[1536] = 0;
        weight_rom[1537] = 1;
        weight_rom[1538] = 2;
        weight_rom[1539] = 2;
        weight_rom[1540] = -3;
        weight_rom[1541] = -2;
        weight_rom[1542] = 0;
        weight_rom[1543] = -3;
        weight_rom[1544] = 3;
        weight_rom[1545] = 31;
        weight_rom[1546] = 47;
        weight_rom[1547] = 3;
        weight_rom[1548] = 37;
        weight_rom[1549] = 30;
        weight_rom[1550] = 45;
        weight_rom[1551] = 6;
        weight_rom[1552] = 27;
        weight_rom[1553] = 92;
        weight_rom[1554] = 59;
        weight_rom[1555] = 49;
        weight_rom[1556] = 66;
        weight_rom[1557] = 98;
        weight_rom[1558] = 75;
        weight_rom[1559] = 50;
        weight_rom[1560] = 10;
        weight_rom[1561] = -20;
        weight_rom[1562] = 2;
        weight_rom[1563] = 0;
        weight_rom[1564] = 3;
        weight_rom[1565] = 1;
        weight_rom[1566] = -3;
        weight_rom[1567] = 2;
        weight_rom[1568] = 2;
        weight_rom[1569] = 1;
        weight_rom[1570] = 2;
        weight_rom[1571] = 0;
        weight_rom[1572] = -1;
        weight_rom[1573] = -1;
        weight_rom[1574] = 3;
        weight_rom[1575] = 1;
        weight_rom[1576] = 2;
        weight_rom[1577] = 0;
        weight_rom[1578] = -3;
        weight_rom[1579] = -1;
        weight_rom[1580] = 2;
        weight_rom[1581] = 6;
        weight_rom[1582] = -18;
        weight_rom[1583] = 0;
        weight_rom[1584] = 0;
        weight_rom[1585] = -3;
        weight_rom[1586] = 0;
        weight_rom[1587] = -3;
        weight_rom[1588] = 0;
        weight_rom[1589] = 0;
        weight_rom[1590] = 0;
        weight_rom[1591] = -2;
        weight_rom[1592] = 2;
        weight_rom[1593] = 2;
        weight_rom[1594] = 3;
        weight_rom[1595] = 2;
        weight_rom[1596] = -2;
        weight_rom[1597] = 1;
        weight_rom[1598] = -2;
        weight_rom[1599] = -3;
        weight_rom[1600] = 2;
        weight_rom[1601] = 3;
        weight_rom[1602] = 28;
        weight_rom[1603] = 40;
        weight_rom[1604] = 38;
        weight_rom[1605] = 42;
        weight_rom[1606] = 51;
        weight_rom[1607] = 60;
        weight_rom[1608] = 83;
        weight_rom[1609] = 65;
        weight_rom[1610] = -9;
        weight_rom[1611] = 12;
        weight_rom[1612] = 48;
        weight_rom[1613] = 48;
        weight_rom[1614] = 54;
        weight_rom[1615] = 36;
        weight_rom[1616] = 34;
        weight_rom[1617] = 31;
        weight_rom[1618] = 38;
        weight_rom[1619] = 25;
        weight_rom[1620] = 1;
        weight_rom[1621] = 2;
        weight_rom[1622] = -2;
        weight_rom[1623] = 0;
        weight_rom[1624] = -2;
        weight_rom[1625] = 1;
        weight_rom[1626] = 1;
        weight_rom[1627] = 3;
        weight_rom[1628] = 24;
        weight_rom[1629] = 3;
        weight_rom[1630] = 40;
        weight_rom[1631] = 70;
        weight_rom[1632] = 75;
        weight_rom[1633] = 75;
        weight_rom[1634] = 103;
        weight_rom[1635] = 98;
        weight_rom[1636] = 78;
        weight_rom[1637] = 28;
        weight_rom[1638] = 33;
        weight_rom[1639] = 2;
        weight_rom[1640] = 55;
        weight_rom[1641] = 63;
        weight_rom[1642] = 115;
        weight_rom[1643] = 67;
        weight_rom[1644] = 71;
        weight_rom[1645] = 54;
        weight_rom[1646] = 48;
        weight_rom[1647] = 40;
        weight_rom[1648] = 14;
        weight_rom[1649] = 2;
        weight_rom[1650] = 0;
        weight_rom[1651] = 3;
        weight_rom[1652] = 2;
        weight_rom[1653] = -3;
        weight_rom[1654] = 21;
        weight_rom[1655] = 0;
        weight_rom[1656] = -2;
        weight_rom[1657] = 28;
        weight_rom[1658] = 51;
        weight_rom[1659] = 74;
        weight_rom[1660] = 104;
        weight_rom[1661] = 97;
        weight_rom[1662] = 88;
        weight_rom[1663] = 112;
        weight_rom[1664] = 109;
        weight_rom[1665] = 104;
        weight_rom[1666] = 91;
        weight_rom[1667] = 80;
        weight_rom[1668] = 59;
        weight_rom[1669] = 68;
        weight_rom[1670] = 79;
        weight_rom[1671] = 62;
        weight_rom[1672] = 81;
        weight_rom[1673] = 38;
        weight_rom[1674] = 18;
        weight_rom[1675] = 53;
        weight_rom[1676] = 65;
        weight_rom[1677] = 22;
        weight_rom[1678] = 0;
        weight_rom[1679] = -3;
        weight_rom[1680] = -2;
        weight_rom[1681] = 2;
        weight_rom[1682] = -21;
        weight_rom[1683] = -2;
        weight_rom[1684] = -1;
        weight_rom[1685] = 7;
        weight_rom[1686] = 19;
        weight_rom[1687] = 41;
        weight_rom[1688] = 29;
        weight_rom[1689] = 49;
        weight_rom[1690] = 61;
        weight_rom[1691] = 42;
        weight_rom[1692] = 37;
        weight_rom[1693] = 25;
        weight_rom[1694] = 31;
        weight_rom[1695] = 30;
        weight_rom[1696] = 17;
        weight_rom[1697] = 28;
        weight_rom[1698] = 34;
        weight_rom[1699] = 9;
        weight_rom[1700] = -17;
        weight_rom[1701] = -13;
        weight_rom[1702] = -25;
        weight_rom[1703] = -1;
        weight_rom[1704] = 0;
        weight_rom[1705] = 25;
        weight_rom[1706] = 7;
        weight_rom[1707] = -1;
        weight_rom[1708] = 2;
        weight_rom[1709] = 3;
        weight_rom[1710] = 0;
        weight_rom[1711] = 19;
        weight_rom[1712] = 10;
        weight_rom[1713] = -37;
        weight_rom[1714] = 9;
        weight_rom[1715] = 9;
        weight_rom[1716] = 12;
        weight_rom[1717] = 19;
        weight_rom[1718] = 42;
        weight_rom[1719] = 21;
        weight_rom[1720] = 17;
        weight_rom[1721] = 17;
        weight_rom[1722] = 17;
        weight_rom[1723] = 26;
        weight_rom[1724] = 32;
        weight_rom[1725] = 31;
        weight_rom[1726] = 22;
        weight_rom[1727] = 3;
        weight_rom[1728] = 17;
        weight_rom[1729] = -6;
        weight_rom[1730] = -8;
        weight_rom[1731] = -2;
        weight_rom[1732] = 6;
        weight_rom[1733] = 35;
        weight_rom[1734] = 19;
        weight_rom[1735] = 2;
        weight_rom[1736] = 2;
        weight_rom[1737] = 3;
        weight_rom[1738] = 25;
        weight_rom[1739] = 39;
        weight_rom[1740] = 6;
        weight_rom[1741] = -5;
        weight_rom[1742] = 11;
        weight_rom[1743] = 15;
        weight_rom[1744] = 13;
        weight_rom[1745] = 17;
        weight_rom[1746] = 11;
        weight_rom[1747] = 9;
        weight_rom[1748] = 17;
        weight_rom[1749] = 18;
        weight_rom[1750] = 14;
        weight_rom[1751] = 17;
        weight_rom[1752] = 16;
        weight_rom[1753] = 8;
        weight_rom[1754] = 12;
        weight_rom[1755] = -2;
        weight_rom[1756] = -8;
        weight_rom[1757] = -3;
        weight_rom[1758] = -10;
        weight_rom[1759] = -3;
        weight_rom[1760] = 36;
        weight_rom[1761] = 34;
        weight_rom[1762] = 19;
        weight_rom[1763] = 24;
        weight_rom[1764] = 1;
        weight_rom[1765] = 34;
        weight_rom[1766] = -11;
        weight_rom[1767] = 25;
        weight_rom[1768] = 14;
        weight_rom[1769] = 26;
        weight_rom[1770] = 16;
        weight_rom[1771] = 10;
        weight_rom[1772] = 17;
        weight_rom[1773] = 10;
        weight_rom[1774] = 9;
        weight_rom[1775] = 12;
        weight_rom[1776] = 11;
        weight_rom[1777] = 6;
        weight_rom[1778] = 21;
        weight_rom[1779] = 11;
        weight_rom[1780] = 2;
        weight_rom[1781] = 11;
        weight_rom[1782] = 3;
        weight_rom[1783] = 2;
        weight_rom[1784] = -14;
        weight_rom[1785] = 2;
        weight_rom[1786] = 3;
        weight_rom[1787] = -6;
        weight_rom[1788] = 29;
        weight_rom[1789] = 44;
        weight_rom[1790] = 15;
        weight_rom[1791] = -5;
        weight_rom[1792] = -13;
        weight_rom[1793] = 7;
        weight_rom[1794] = 12;
        weight_rom[1795] = 7;
        weight_rom[1796] = 12;
        weight_rom[1797] = 16;
        weight_rom[1798] = 11;
        weight_rom[1799] = 7;
        weight_rom[1800] = -3;
        weight_rom[1801] = 9;
        weight_rom[1802] = 12;
        weight_rom[1803] = 11;
        weight_rom[1804] = 3;
        weight_rom[1805] = 7;
        weight_rom[1806] = 11;
        weight_rom[1807] = 10;
        weight_rom[1808] = 15;
        weight_rom[1809] = 14;
        weight_rom[1810] = -1;
        weight_rom[1811] = 14;
        weight_rom[1812] = 21;
        weight_rom[1813] = 0;
        weight_rom[1814] = 12;
        weight_rom[1815] = 12;
        weight_rom[1816] = 27;
        weight_rom[1817] = 26;
        weight_rom[1818] = 20;
        weight_rom[1819] = 12;
        weight_rom[1820] = -1;
        weight_rom[1821] = 12;
        weight_rom[1822] = 23;
        weight_rom[1823] = 9;
        weight_rom[1824] = 8;
        weight_rom[1825] = 12;
        weight_rom[1826] = -9;
        weight_rom[1827] = 0;
        weight_rom[1828] = 1;
        weight_rom[1829] = -3;
        weight_rom[1830] = -11;
        weight_rom[1831] = -11;
        weight_rom[1832] = -17;
        weight_rom[1833] = -8;
        weight_rom[1834] = 6;
        weight_rom[1835] = -4;
        weight_rom[1836] = -5;
        weight_rom[1837] = -7;
        weight_rom[1838] = 7;
        weight_rom[1839] = 7;
        weight_rom[1840] = 12;
        weight_rom[1841] = 9;
        weight_rom[1842] = 25;
        weight_rom[1843] = 6;
        weight_rom[1844] = 45;
        weight_rom[1845] = 54;
        weight_rom[1846] = -3;
        weight_rom[1847] = -26;
        weight_rom[1848] = -9;
        weight_rom[1849] = -29;
        weight_rom[1850] = 21;
        weight_rom[1851] = 35;
        weight_rom[1852] = 4;
        weight_rom[1853] = 10;
        weight_rom[1854] = -3;
        weight_rom[1855] = -12;
        weight_rom[1856] = -28;
        weight_rom[1857] = -17;
        weight_rom[1858] = -27;
        weight_rom[1859] = -23;
        weight_rom[1860] = -31;
        weight_rom[1861] = -15;
        weight_rom[1862] = -13;
        weight_rom[1863] = -22;
        weight_rom[1864] = -2;
        weight_rom[1865] = 4;
        weight_rom[1866] = 6;
        weight_rom[1867] = -1;
        weight_rom[1868] = 19;
        weight_rom[1869] = 4;
        weight_rom[1870] = 1;
        weight_rom[1871] = 27;
        weight_rom[1872] = 74;
        weight_rom[1873] = 64;
        weight_rom[1874] = 48;
        weight_rom[1875] = 19;
        weight_rom[1876] = -28;
        weight_rom[1877] = -7;
        weight_rom[1878] = 22;
        weight_rom[1879] = 22;
        weight_rom[1880] = 12;
        weight_rom[1881] = -14;
        weight_rom[1882] = -15;
        weight_rom[1883] = -26;
        weight_rom[1884] = -24;
        weight_rom[1885] = -29;
        weight_rom[1886] = -32;
        weight_rom[1887] = -21;
        weight_rom[1888] = -24;
        weight_rom[1889] = -20;
        weight_rom[1890] = -30;
        weight_rom[1891] = -52;
        weight_rom[1892] = -31;
        weight_rom[1893] = -5;
        weight_rom[1894] = 1;
        weight_rom[1895] = 16;
        weight_rom[1896] = 0;
        weight_rom[1897] = -8;
        weight_rom[1898] = -21;
        weight_rom[1899] = 16;
        weight_rom[1900] = 30;
        weight_rom[1901] = 40;
        weight_rom[1902] = 13;
        weight_rom[1903] = -5;
        weight_rom[1904] = -14;
        weight_rom[1905] = -4;
        weight_rom[1906] = 2;
        weight_rom[1907] = 18;
        weight_rom[1908] = -11;
        weight_rom[1909] = -26;
        weight_rom[1910] = -29;
        weight_rom[1911] = -21;
        weight_rom[1912] = -22;
        weight_rom[1913] = -14;
        weight_rom[1914] = 10;
        weight_rom[1915] = 2;
        weight_rom[1916] = 3;
        weight_rom[1917] = -5;
        weight_rom[1918] = -31;
        weight_rom[1919] = -28;
        weight_rom[1920] = -23;
        weight_rom[1921] = -6;
        weight_rom[1922] = -5;
        weight_rom[1923] = -7;
        weight_rom[1924] = -12;
        weight_rom[1925] = -27;
        weight_rom[1926] = -40;
        weight_rom[1927] = -11;
        weight_rom[1928] = 39;
        weight_rom[1929] = 19;
        weight_rom[1930] = 28;
        weight_rom[1931] = -3;
        weight_rom[1932] = -2;
        weight_rom[1933] = -5;
        weight_rom[1934] = 7;
        weight_rom[1935] = 26;
        weight_rom[1936] = -46;
        weight_rom[1937] = -29;
        weight_rom[1938] = -8;
        weight_rom[1939] = -22;
        weight_rom[1940] = -3;
        weight_rom[1941] = 4;
        weight_rom[1942] = 19;
        weight_rom[1943] = 27;
        weight_rom[1944] = 17;
        weight_rom[1945] = 13;
        weight_rom[1946] = -12;
        weight_rom[1947] = -37;
        weight_rom[1948] = -28;
        weight_rom[1949] = -10;
        weight_rom[1950] = -1;
        weight_rom[1951] = 6;
        weight_rom[1952] = -31;
        weight_rom[1953] = -30;
        weight_rom[1954] = -13;
        weight_rom[1955] = 37;
        weight_rom[1956] = 44;
        weight_rom[1957] = 25;
        weight_rom[1958] = -10;
        weight_rom[1959] = 10;
        weight_rom[1960] = -3;
        weight_rom[1961] = 6;
        weight_rom[1962] = -16;
        weight_rom[1963] = -9;
        weight_rom[1964] = -61;
        weight_rom[1965] = -10;
        weight_rom[1966] = -5;
        weight_rom[1967] = 1;
        weight_rom[1968] = 15;
        weight_rom[1969] = 18;
        weight_rom[1970] = 27;
        weight_rom[1971] = 17;
        weight_rom[1972] = 14;
        weight_rom[1973] = 7;
        weight_rom[1974] = -11;
        weight_rom[1975] = -12;
        weight_rom[1976] = -22;
        weight_rom[1977] = -11;
        weight_rom[1978] = -3;
        weight_rom[1979] = -19;
        weight_rom[1980] = -7;
        weight_rom[1981] = 9;
        weight_rom[1982] = 7;
        weight_rom[1983] = 30;
        weight_rom[1984] = 70;
        weight_rom[1985] = -2;
        weight_rom[1986] = 16;
        weight_rom[1987] = 2;
        weight_rom[1988] = 0;
        weight_rom[1989] = 21;
        weight_rom[1990] = 17;
        weight_rom[1991] = -19;
        weight_rom[1992] = -19;
        weight_rom[1993] = 11;
        weight_rom[1994] = -8;
        weight_rom[1995] = 10;
        weight_rom[1996] = 2;
        weight_rom[1997] = 16;
        weight_rom[1998] = 22;
        weight_rom[1999] = 13;
        weight_rom[2000] = 9;
        weight_rom[2001] = 0;
        weight_rom[2002] = -8;
        weight_rom[2003] = -19;
        weight_rom[2004] = -18;
        weight_rom[2005] = -7;
        weight_rom[2006] = -7;
        weight_rom[2007] = 9;
        weight_rom[2008] = 14;
        weight_rom[2009] = 16;
        weight_rom[2010] = 11;
        weight_rom[2011] = 42;
        weight_rom[2012] = 70;
        weight_rom[2013] = 34;
        weight_rom[2014] = -24;
        weight_rom[2015] = 13;
        weight_rom[2016] = -2;
        weight_rom[2017] = 0;
        weight_rom[2018] = 59;
        weight_rom[2019] = 25;
        weight_rom[2020] = 16;
        weight_rom[2021] = 0;
        weight_rom[2022] = -11;
        weight_rom[2023] = -5;
        weight_rom[2024] = -14;
        weight_rom[2025] = 12;
        weight_rom[2026] = 2;
        weight_rom[2027] = 17;
        weight_rom[2028] = 8;
        weight_rom[2029] = 7;
        weight_rom[2030] = -9;
        weight_rom[2031] = -20;
        weight_rom[2032] = -22;
        weight_rom[2033] = 6;
        weight_rom[2034] = 19;
        weight_rom[2035] = 30;
        weight_rom[2036] = 19;
        weight_rom[2037] = 32;
        weight_rom[2038] = 31;
        weight_rom[2039] = 24;
        weight_rom[2040] = 56;
        weight_rom[2041] = 28;
        weight_rom[2042] = -26;
        weight_rom[2043] = -36;
        weight_rom[2044] = -2;
        weight_rom[2045] = 4;
        weight_rom[2046] = -2;
        weight_rom[2047] = 52;
        weight_rom[2048] = 33;
        weight_rom[2049] = 22;
        weight_rom[2050] = 28;
        weight_rom[2051] = 8;
        weight_rom[2052] = -11;
        weight_rom[2053] = -18;
        weight_rom[2054] = 5;
        weight_rom[2055] = 0;
        weight_rom[2056] = -16;
        weight_rom[2057] = -32;
        weight_rom[2058] = -36;
        weight_rom[2059] = -15;
        weight_rom[2060] = 6;
        weight_rom[2061] = 26;
        weight_rom[2062] = 31;
        weight_rom[2063] = 29;
        weight_rom[2064] = 20;
        weight_rom[2065] = 9;
        weight_rom[2066] = 23;
        weight_rom[2067] = 23;
        weight_rom[2068] = 12;
        weight_rom[2069] = 35;
        weight_rom[2070] = 39;
        weight_rom[2071] = 0;
        weight_rom[2072] = -2;
        weight_rom[2073] = 3;
        weight_rom[2074] = 39;
        weight_rom[2075] = 39;
        weight_rom[2076] = 18;
        weight_rom[2077] = 27;
        weight_rom[2078] = 32;
        weight_rom[2079] = 26;
        weight_rom[2080] = 10;
        weight_rom[2081] = -6;
        weight_rom[2082] = 1;
        weight_rom[2083] = -7;
        weight_rom[2084] = -12;
        weight_rom[2085] = -23;
        weight_rom[2086] = -28;
        weight_rom[2087] = 3;
        weight_rom[2088] = 31;
        weight_rom[2089] = 40;
        weight_rom[2090] = 24;
        weight_rom[2091] = 30;
        weight_rom[2092] = 0;
        weight_rom[2093] = 10;
        weight_rom[2094] = 49;
        weight_rom[2095] = 36;
        weight_rom[2096] = 49;
        weight_rom[2097] = 76;
        weight_rom[2098] = -6;
        weight_rom[2099] = -35;
        weight_rom[2100] = -3;
        weight_rom[2101] = 2;
        weight_rom[2102] = -7;
        weight_rom[2103] = 49;
        weight_rom[2104] = 50;
        weight_rom[2105] = 31;
        weight_rom[2106] = 37;
        weight_rom[2107] = 37;
        weight_rom[2108] = 25;
        weight_rom[2109] = 19;
        weight_rom[2110] = 21;
        weight_rom[2111] = 15;
        weight_rom[2112] = 23;
        weight_rom[2113] = 11;
        weight_rom[2114] = 5;
        weight_rom[2115] = 24;
        weight_rom[2116] = 26;
        weight_rom[2117] = 31;
        weight_rom[2118] = 32;
        weight_rom[2119] = 19;
        weight_rom[2120] = 26;
        weight_rom[2121] = 33;
        weight_rom[2122] = 38;
        weight_rom[2123] = 29;
        weight_rom[2124] = 36;
        weight_rom[2125] = 34;
        weight_rom[2126] = 8;
        weight_rom[2127] = -18;
        weight_rom[2128] = 2;
        weight_rom[2129] = 33;
        weight_rom[2130] = -6;
        weight_rom[2131] = 61;
        weight_rom[2132] = 55;
        weight_rom[2133] = 59;
        weight_rom[2134] = 32;
        weight_rom[2135] = 25;
        weight_rom[2136] = 37;
        weight_rom[2137] = 33;
        weight_rom[2138] = 28;
        weight_rom[2139] = 14;
        weight_rom[2140] = 13;
        weight_rom[2141] = 12;
        weight_rom[2142] = 12;
        weight_rom[2143] = 15;
        weight_rom[2144] = 17;
        weight_rom[2145] = 18;
        weight_rom[2146] = 26;
        weight_rom[2147] = 20;
        weight_rom[2148] = 27;
        weight_rom[2149] = 34;
        weight_rom[2150] = 34;
        weight_rom[2151] = 37;
        weight_rom[2152] = 14;
        weight_rom[2153] = 16;
        weight_rom[2154] = 10;
        weight_rom[2155] = 0;
        weight_rom[2156] = 3;
        weight_rom[2157] = 11;
        weight_rom[2158] = 31;
        weight_rom[2159] = 72;
        weight_rom[2160] = 48;
        weight_rom[2161] = 20;
        weight_rom[2162] = 7;
        weight_rom[2163] = 27;
        weight_rom[2164] = 16;
        weight_rom[2165] = 4;
        weight_rom[2166] = 10;
        weight_rom[2167] = 17;
        weight_rom[2168] = 16;
        weight_rom[2169] = 29;
        weight_rom[2170] = 18;
        weight_rom[2171] = 22;
        weight_rom[2172] = 13;
        weight_rom[2173] = 19;
        weight_rom[2174] = 26;
        weight_rom[2175] = 20;
        weight_rom[2176] = 9;
        weight_rom[2177] = 13;
        weight_rom[2178] = 38;
        weight_rom[2179] = 48;
        weight_rom[2180] = -22;
        weight_rom[2181] = 3;
        weight_rom[2182] = 37;
        weight_rom[2183] = 2;
        weight_rom[2184] = 0;
        weight_rom[2185] = -3;
        weight_rom[2186] = 54;
        weight_rom[2187] = 75;
        weight_rom[2188] = 28;
        weight_rom[2189] = -20;
        weight_rom[2190] = 3;
        weight_rom[2191] = 4;
        weight_rom[2192] = 7;
        weight_rom[2193] = 16;
        weight_rom[2194] = 5;
        weight_rom[2195] = 20;
        weight_rom[2196] = 24;
        weight_rom[2197] = 26;
        weight_rom[2198] = 10;
        weight_rom[2199] = 23;
        weight_rom[2200] = 14;
        weight_rom[2201] = 4;
        weight_rom[2202] = 16;
        weight_rom[2203] = 22;
        weight_rom[2204] = 22;
        weight_rom[2205] = 17;
        weight_rom[2206] = 29;
        weight_rom[2207] = -3;
        weight_rom[2208] = -26;
        weight_rom[2209] = 0;
        weight_rom[2210] = -3;
        weight_rom[2211] = -3;
        weight_rom[2212] = -2;
        weight_rom[2213] = -2;
        weight_rom[2214] = 34;
        weight_rom[2215] = 77;
        weight_rom[2216] = 27;
        weight_rom[2217] = 16;
        weight_rom[2218] = 11;
        weight_rom[2219] = 15;
        weight_rom[2220] = 14;
        weight_rom[2221] = 24;
        weight_rom[2222] = 32;
        weight_rom[2223] = 26;
        weight_rom[2224] = 17;
        weight_rom[2225] = 14;
        weight_rom[2226] = 20;
        weight_rom[2227] = 13;
        weight_rom[2228] = -1;
        weight_rom[2229] = 1;
        weight_rom[2230] = 16;
        weight_rom[2231] = 14;
        weight_rom[2232] = 16;
        weight_rom[2233] = 4;
        weight_rom[2234] = 9;
        weight_rom[2235] = 20;
        weight_rom[2236] = 4;
        weight_rom[2237] = 30;
        weight_rom[2238] = -25;
        weight_rom[2239] = 1;
        weight_rom[2240] = -1;
        weight_rom[2241] = 3;
        weight_rom[2242] = 18;
        weight_rom[2243] = 50;
        weight_rom[2244] = 52;
        weight_rom[2245] = 4;
        weight_rom[2246] = 18;
        weight_rom[2247] = 24;
        weight_rom[2248] = 2;
        weight_rom[2249] = 25;
        weight_rom[2250] = 18;
        weight_rom[2251] = 33;
        weight_rom[2252] = 33;
        weight_rom[2253] = 43;
        weight_rom[2254] = 38;
        weight_rom[2255] = 24;
        weight_rom[2256] = 25;
        weight_rom[2257] = 27;
        weight_rom[2258] = 4;
        weight_rom[2259] = -10;
        weight_rom[2260] = -22;
        weight_rom[2261] = 0;
        weight_rom[2262] = -13;
        weight_rom[2263] = -28;
        weight_rom[2264] = 20;
        weight_rom[2265] = 32;
        weight_rom[2266] = 3;
        weight_rom[2267] = 0;
        weight_rom[2268] = 3;
        weight_rom[2269] = -1;
        weight_rom[2270] = 1;
        weight_rom[2271] = -6;
        weight_rom[2272] = 11;
        weight_rom[2273] = 1;
        weight_rom[2274] = 37;
        weight_rom[2275] = 6;
        weight_rom[2276] = 32;
        weight_rom[2277] = 11;
        weight_rom[2278] = 23;
        weight_rom[2279] = 13;
        weight_rom[2280] = 25;
        weight_rom[2281] = 21;
        weight_rom[2282] = 3;
        weight_rom[2283] = 18;
        weight_rom[2284] = 4;
        weight_rom[2285] = 2;
        weight_rom[2286] = -23;
        weight_rom[2287] = -6;
        weight_rom[2288] = -58;
        weight_rom[2289] = -46;
        weight_rom[2290] = -1;
        weight_rom[2291] = -4;
        weight_rom[2292] = 15;
        weight_rom[2293] = -2;
        weight_rom[2294] = -2;
        weight_rom[2295] = 2;
        weight_rom[2296] = 1;
        weight_rom[2297] = 3;
        weight_rom[2298] = 1;
        weight_rom[2299] = -1;
        weight_rom[2300] = -30;
        weight_rom[2301] = -50;
        weight_rom[2302] = -17;
        weight_rom[2303] = -13;
        weight_rom[2304] = -18;
        weight_rom[2305] = 1;
        weight_rom[2306] = -11;
        weight_rom[2307] = -6;
        weight_rom[2308] = 10;
        weight_rom[2309] = 13;
        weight_rom[2310] = -12;
        weight_rom[2311] = 17;
        weight_rom[2312] = 15;
        weight_rom[2313] = -6;
        weight_rom[2314] = -17;
        weight_rom[2315] = -12;
        weight_rom[2316] = -21;
        weight_rom[2317] = -3;
        weight_rom[2318] = -23;
        weight_rom[2319] = -12;
        weight_rom[2320] = -2;
        weight_rom[2321] = 3;
        weight_rom[2322] = -1;
        weight_rom[2323] = 0;
        weight_rom[2324] = -3;
        weight_rom[2325] = 0;
        weight_rom[2326] = -3;
        weight_rom[2327] = 2;
        weight_rom[2328] = -2;
        weight_rom[2329] = -5;
        weight_rom[2330] = -1;
        weight_rom[2331] = 1;
        weight_rom[2332] = 5;
        weight_rom[2333] = -1;
        weight_rom[2334] = -12;
        weight_rom[2335] = 35;
        weight_rom[2336] = 28;
        weight_rom[2337] = 5;
        weight_rom[2338] = -21;
        weight_rom[2339] = -17;
        weight_rom[2340] = 3;
        weight_rom[2341] = 13;
        weight_rom[2342] = -7;
        weight_rom[2343] = 0;
        weight_rom[2344] = -17;
        weight_rom[2345] = -3;
        weight_rom[2346] = -28;
        weight_rom[2347] = 2;
        weight_rom[2348] = -2;
        weight_rom[2349] = -3;
        weight_rom[2350] = 2;
        weight_rom[2351] = 1;
        weight_rom[2352] = 0;
        weight_rom[2353] = -2;
        weight_rom[2354] = 2;
        weight_rom[2355] = -3;
        weight_rom[2356] = -1;
        weight_rom[2357] = -2;
        weight_rom[2358] = 3;
        weight_rom[2359] = -3;
        weight_rom[2360] = 3;
        weight_rom[2361] = -3;
        weight_rom[2362] = -1;
        weight_rom[2363] = 3;
        weight_rom[2364] = -2;
        weight_rom[2365] = -24;
        weight_rom[2366] = -21;
        weight_rom[2367] = -1;
        weight_rom[2368] = -1;
        weight_rom[2369] = 0;
        weight_rom[2370] = 3;
        weight_rom[2371] = -3;
        weight_rom[2372] = 2;
        weight_rom[2373] = -1;
        weight_rom[2374] = 0;
        weight_rom[2375] = 1;
        weight_rom[2376] = 0;
        weight_rom[2377] = 2;
        weight_rom[2378] = -1;
        weight_rom[2379] = 2;
        weight_rom[2380] = -2;
        weight_rom[2381] = 3;
        weight_rom[2382] = -3;
        weight_rom[2383] = 0;
        weight_rom[2384] = -2;
        weight_rom[2385] = 0;
        weight_rom[2386] = -16;
        weight_rom[2387] = -36;
        weight_rom[2388] = -21;
        weight_rom[2389] = -8;
        weight_rom[2390] = -30;
        weight_rom[2391] = -23;
        weight_rom[2392] = -49;
        weight_rom[2393] = -31;
        weight_rom[2394] = 1;
        weight_rom[2395] = -22;
        weight_rom[2396] = -56;
        weight_rom[2397] = -20;
        weight_rom[2398] = -5;
        weight_rom[2399] = -23;
        weight_rom[2400] = -18;
        weight_rom[2401] = -28;
        weight_rom[2402] = -41;
        weight_rom[2403] = -25;
        weight_rom[2404] = 2;
        weight_rom[2405] = 2;
        weight_rom[2406] = -2;
        weight_rom[2407] = 1;
        weight_rom[2408] = -1;
        weight_rom[2409] = -1;
        weight_rom[2410] = 2;
        weight_rom[2411] = -3;
        weight_rom[2412] = 10;
        weight_rom[2413] = -1;
        weight_rom[2414] = -1;
        weight_rom[2415] = -34;
        weight_rom[2416] = -45;
        weight_rom[2417] = -47;
        weight_rom[2418] = -59;
        weight_rom[2419] = -42;
        weight_rom[2420] = -36;
        weight_rom[2421] = -12;
        weight_rom[2422] = -18;
        weight_rom[2423] = -30;
        weight_rom[2424] = -23;
        weight_rom[2425] = -18;
        weight_rom[2426] = -5;
        weight_rom[2427] = 15;
        weight_rom[2428] = 3;
        weight_rom[2429] = -2;
        weight_rom[2430] = -8;
        weight_rom[2431] = -26;
        weight_rom[2432] = -20;
        weight_rom[2433] = -23;
        weight_rom[2434] = 0;
        weight_rom[2435] = 0;
        weight_rom[2436] = 2;
        weight_rom[2437] = -3;
        weight_rom[2438] = -17;
        weight_rom[2439] = 1;
        weight_rom[2440] = -1;
        weight_rom[2441] = 22;
        weight_rom[2442] = 6;
        weight_rom[2443] = -9;
        weight_rom[2444] = -10;
        weight_rom[2445] = -42;
        weight_rom[2446] = -7;
        weight_rom[2447] = -17;
        weight_rom[2448] = -12;
        weight_rom[2449] = -33;
        weight_rom[2450] = -12;
        weight_rom[2451] = -13;
        weight_rom[2452] = -9;
        weight_rom[2453] = 6;
        weight_rom[2454] = 24;
        weight_rom[2455] = 30;
        weight_rom[2456] = 31;
        weight_rom[2457] = 23;
        weight_rom[2458] = 6;
        weight_rom[2459] = 19;
        weight_rom[2460] = 7;
        weight_rom[2461] = -5;
        weight_rom[2462] = 0;
        weight_rom[2463] = 0;
        weight_rom[2464] = 2;
        weight_rom[2465] = 0;
        weight_rom[2466] = -6;
        weight_rom[2467] = 2;
        weight_rom[2468] = 40;
        weight_rom[2469] = 40;
        weight_rom[2470] = -1;
        weight_rom[2471] = 15;
        weight_rom[2472] = 5;
        weight_rom[2473] = -4;
        weight_rom[2474] = 7;
        weight_rom[2475] = 14;
        weight_rom[2476] = 11;
        weight_rom[2477] = 1;
        weight_rom[2478] = -3;
        weight_rom[2479] = -10;
        weight_rom[2480] = 10;
        weight_rom[2481] = -3;
        weight_rom[2482] = 3;
        weight_rom[2483] = 7;
        weight_rom[2484] = -3;
        weight_rom[2485] = 8;
        weight_rom[2486] = 18;
        weight_rom[2487] = 29;
        weight_rom[2488] = 86;
        weight_rom[2489] = 24;
        weight_rom[2490] = 29;
        weight_rom[2491] = 0;
        weight_rom[2492] = 0;
        weight_rom[2493] = 3;
        weight_rom[2494] = -3;
        weight_rom[2495] = 25;
        weight_rom[2496] = 18;
        weight_rom[2497] = 44;
        weight_rom[2498] = 23;
        weight_rom[2499] = 26;
        weight_rom[2500] = 14;
        weight_rom[2501] = 23;
        weight_rom[2502] = 9;
        weight_rom[2503] = 24;
        weight_rom[2504] = 20;
        weight_rom[2505] = 15;
        weight_rom[2506] = 8;
        weight_rom[2507] = 10;
        weight_rom[2508] = 7;
        weight_rom[2509] = 2;
        weight_rom[2510] = -10;
        weight_rom[2511] = 6;
        weight_rom[2512] = -12;
        weight_rom[2513] = -20;
        weight_rom[2514] = -3;
        weight_rom[2515] = 25;
        weight_rom[2516] = 29;
        weight_rom[2517] = 57;
        weight_rom[2518] = 43;
        weight_rom[2519] = 0;
        weight_rom[2520] = 1;
        weight_rom[2521] = 0;
        weight_rom[2522] = 27;
        weight_rom[2523] = 23;
        weight_rom[2524] = 43;
        weight_rom[2525] = 19;
        weight_rom[2526] = 28;
        weight_rom[2527] = 4;
        weight_rom[2528] = 23;
        weight_rom[2529] = 17;
        weight_rom[2530] = 25;
        weight_rom[2531] = 20;
        weight_rom[2532] = 7;
        weight_rom[2533] = 14;
        weight_rom[2534] = 15;
        weight_rom[2535] = 26;
        weight_rom[2536] = 12;
        weight_rom[2537] = 4;
        weight_rom[2538] = -2;
        weight_rom[2539] = 0;
        weight_rom[2540] = 1;
        weight_rom[2541] = -9;
        weight_rom[2542] = -6;
        weight_rom[2543] = 6;
        weight_rom[2544] = 48;
        weight_rom[2545] = 98;
        weight_rom[2546] = 47;
        weight_rom[2547] = -25;
        weight_rom[2548] = -2;
        weight_rom[2549] = 34;
        weight_rom[2550] = -24;
        weight_rom[2551] = 30;
        weight_rom[2552] = 11;
        weight_rom[2553] = 24;
        weight_rom[2554] = 10;
        weight_rom[2555] = 17;
        weight_rom[2556] = 11;
        weight_rom[2557] = 14;
        weight_rom[2558] = 6;
        weight_rom[2559] = 0;
        weight_rom[2560] = 14;
        weight_rom[2561] = 10;
        weight_rom[2562] = 19;
        weight_rom[2563] = 27;
        weight_rom[2564] = 19;
        weight_rom[2565] = 20;
        weight_rom[2566] = 4;
        weight_rom[2567] = 7;
        weight_rom[2568] = 2;
        weight_rom[2569] = -5;
        weight_rom[2570] = -15;
        weight_rom[2571] = 4;
        weight_rom[2572] = 29;
        weight_rom[2573] = 83;
        weight_rom[2574] = 41;
        weight_rom[2575] = 2;
        weight_rom[2576] = -6;
        weight_rom[2577] = 12;
        weight_rom[2578] = 12;
        weight_rom[2579] = 11;
        weight_rom[2580] = 24;
        weight_rom[2581] = 22;
        weight_rom[2582] = 15;
        weight_rom[2583] = 7;
        weight_rom[2584] = 5;
        weight_rom[2585] = 1;
        weight_rom[2586] = -6;
        weight_rom[2587] = 3;
        weight_rom[2588] = -2;
        weight_rom[2589] = 4;
        weight_rom[2590] = 4;
        weight_rom[2591] = -5;
        weight_rom[2592] = 5;
        weight_rom[2593] = 10;
        weight_rom[2594] = 17;
        weight_rom[2595] = 8;
        weight_rom[2596] = 10;
        weight_rom[2597] = 13;
        weight_rom[2598] = 7;
        weight_rom[2599] = -15;
        weight_rom[2600] = 48;
        weight_rom[2601] = 99;
        weight_rom[2602] = 53;
        weight_rom[2603] = 21;
        weight_rom[2604] = -2;
        weight_rom[2605] = 15;
        weight_rom[2606] = 12;
        weight_rom[2607] = 19;
        weight_rom[2608] = 30;
        weight_rom[2609] = 7;
        weight_rom[2610] = 16;
        weight_rom[2611] = 8;
        weight_rom[2612] = 1;
        weight_rom[2613] = 3;
        weight_rom[2614] = -12;
        weight_rom[2615] = -13;
        weight_rom[2616] = -9;
        weight_rom[2617] = -16;
        weight_rom[2618] = -8;
        weight_rom[2619] = 10;
        weight_rom[2620] = -4;
        weight_rom[2621] = 8;
        weight_rom[2622] = 7;
        weight_rom[2623] = 16;
        weight_rom[2624] = 21;
        weight_rom[2625] = 23;
        weight_rom[2626] = 25;
        weight_rom[2627] = 5;
        weight_rom[2628] = 11;
        weight_rom[2629] = 96;
        weight_rom[2630] = 57;
        weight_rom[2631] = 25;
        weight_rom[2632] = -4;
        weight_rom[2633] = -2;
        weight_rom[2634] = -22;
        weight_rom[2635] = 26;
        weight_rom[2636] = 1;
        weight_rom[2637] = -15;
        weight_rom[2638] = -11;
        weight_rom[2639] = 9;
        weight_rom[2640] = -12;
        weight_rom[2641] = -18;
        weight_rom[2642] = -19;
        weight_rom[2643] = -29;
        weight_rom[2644] = -33;
        weight_rom[2645] = -16;
        weight_rom[2646] = -21;
        weight_rom[2647] = -12;
        weight_rom[2648] = 10;
        weight_rom[2649] = 4;
        weight_rom[2650] = 9;
        weight_rom[2651] = 14;
        weight_rom[2652] = 8;
        weight_rom[2653] = 14;
        weight_rom[2654] = -4;
        weight_rom[2655] = 4;
        weight_rom[2656] = -19;
        weight_rom[2657] = 60;
        weight_rom[2658] = 35;
        weight_rom[2659] = -6;
        weight_rom[2660] = -3;
        weight_rom[2661] = -17;
        weight_rom[2662] = -9;
        weight_rom[2663] = 28;
        weight_rom[2664] = 13;
        weight_rom[2665] = 0;
        weight_rom[2666] = -3;
        weight_rom[2667] = -11;
        weight_rom[2668] = -12;
        weight_rom[2669] = 2;
        weight_rom[2670] = 15;
        weight_rom[2671] = 5;
        weight_rom[2672] = 15;
        weight_rom[2673] = -17;
        weight_rom[2674] = -4;
        weight_rom[2675] = 18;
        weight_rom[2676] = 21;
        weight_rom[2677] = 39;
        weight_rom[2678] = 26;
        weight_rom[2679] = 20;
        weight_rom[2680] = 11;
        weight_rom[2681] = -7;
        weight_rom[2682] = 0;
        weight_rom[2683] = -24;
        weight_rom[2684] = -12;
        weight_rom[2685] = 36;
        weight_rom[2686] = 79;
        weight_rom[2687] = 13;
        weight_rom[2688] = 1;
        weight_rom[2689] = 2;
        weight_rom[2690] = -13;
        weight_rom[2691] = 2;
        weight_rom[2692] = 21;
        weight_rom[2693] = 12;
        weight_rom[2694] = 12;
        weight_rom[2695] = 19;
        weight_rom[2696] = 14;
        weight_rom[2697] = 13;
        weight_rom[2698] = 23;
        weight_rom[2699] = 25;
        weight_rom[2700] = 14;
        weight_rom[2701] = 1;
        weight_rom[2702] = 15;
        weight_rom[2703] = 30;
        weight_rom[2704] = 39;
        weight_rom[2705] = 34;
        weight_rom[2706] = 30;
        weight_rom[2707] = 17;
        weight_rom[2708] = 1;
        weight_rom[2709] = -10;
        weight_rom[2710] = -25;
        weight_rom[2711] = -12;
        weight_rom[2712] = -54;
        weight_rom[2713] = -18;
        weight_rom[2714] = -13;
        weight_rom[2715] = 13;
        weight_rom[2716] = -2;
        weight_rom[2717] = -7;
        weight_rom[2718] = -26;
        weight_rom[2719] = 0;
        weight_rom[2720] = 53;
        weight_rom[2721] = 34;
        weight_rom[2722] = 17;
        weight_rom[2723] = 30;
        weight_rom[2724] = 17;
        weight_rom[2725] = 27;
        weight_rom[2726] = 21;
        weight_rom[2727] = 15;
        weight_rom[2728] = 10;
        weight_rom[2729] = 25;
        weight_rom[2730] = 22;
        weight_rom[2731] = 34;
        weight_rom[2732] = 41;
        weight_rom[2733] = 32;
        weight_rom[2734] = 31;
        weight_rom[2735] = 13;
        weight_rom[2736] = 2;
        weight_rom[2737] = 3;
        weight_rom[2738] = -11;
        weight_rom[2739] = -36;
        weight_rom[2740] = -26;
        weight_rom[2741] = -57;
        weight_rom[2742] = -29;
        weight_rom[2743] = -25;
        weight_rom[2744] = 2;
        weight_rom[2745] = -11;
        weight_rom[2746] = -5;
        weight_rom[2747] = 27;
        weight_rom[2748] = 41;
        weight_rom[2749] = -2;
        weight_rom[2750] = 6;
        weight_rom[2751] = -8;
        weight_rom[2752] = 14;
        weight_rom[2753] = 15;
        weight_rom[2754] = 15;
        weight_rom[2755] = 9;
        weight_rom[2756] = 17;
        weight_rom[2757] = 9;
        weight_rom[2758] = 16;
        weight_rom[2759] = 12;
        weight_rom[2760] = 24;
        weight_rom[2761] = 35;
        weight_rom[2762] = 25;
        weight_rom[2763] = 21;
        weight_rom[2764] = 8;
        weight_rom[2765] = -3;
        weight_rom[2766] = -13;
        weight_rom[2767] = -13;
        weight_rom[2768] = -29;
        weight_rom[2769] = -23;
        weight_rom[2770] = -63;
        weight_rom[2771] = -1;
        weight_rom[2772] = 0;
        weight_rom[2773] = 26;
        weight_rom[2774] = 29;
        weight_rom[2775] = 2;
        weight_rom[2776] = -10;
        weight_rom[2777] = -23;
        weight_rom[2778] = 6;
        weight_rom[2779] = -10;
        weight_rom[2780] = -14;
        weight_rom[2781] = -5;
        weight_rom[2782] = 2;
        weight_rom[2783] = 11;
        weight_rom[2784] = 26;
        weight_rom[2785] = 13;
        weight_rom[2786] = 4;
        weight_rom[2787] = 24;
        weight_rom[2788] = 27;
        weight_rom[2789] = 29;
        weight_rom[2790] = 24;
        weight_rom[2791] = 20;
        weight_rom[2792] = 21;
        weight_rom[2793] = 10;
        weight_rom[2794] = 17;
        weight_rom[2795] = 15;
        weight_rom[2796] = -31;
        weight_rom[2797] = -54;
        weight_rom[2798] = -34;
        weight_rom[2799] = -17;
        weight_rom[2800] = -2;
        weight_rom[2801] = 0;
        weight_rom[2802] = 38;
        weight_rom[2803] = -21;
        weight_rom[2804] = -7;
        weight_rom[2805] = -13;
        weight_rom[2806] = -5;
        weight_rom[2807] = -10;
        weight_rom[2808] = -10;
        weight_rom[2809] = -5;
        weight_rom[2810] = -11;
        weight_rom[2811] = 3;
        weight_rom[2812] = 24;
        weight_rom[2813] = 18;
        weight_rom[2814] = -12;
        weight_rom[2815] = 9;
        weight_rom[2816] = 22;
        weight_rom[2817] = 21;
        weight_rom[2818] = 18;
        weight_rom[2819] = 21;
        weight_rom[2820] = 1;
        weight_rom[2821] = -16;
        weight_rom[2822] = 7;
        weight_rom[2823] = 19;
        weight_rom[2824] = 2;
        weight_rom[2825] = -68;
        weight_rom[2826] = -64;
        weight_rom[2827] = -35;
        weight_rom[2828] = -2;
        weight_rom[2829] = 7;
        weight_rom[2830] = -9;
        weight_rom[2831] = -2;
        weight_rom[2832] = 6;
        weight_rom[2833] = -5;
        weight_rom[2834] = -11;
        weight_rom[2835] = 6;
        weight_rom[2836] = 4;
        weight_rom[2837] = -17;
        weight_rom[2838] = -28;
        weight_rom[2839] = -16;
        weight_rom[2840] = -3;
        weight_rom[2841] = -7;
        weight_rom[2842] = -1;
        weight_rom[2843] = 9;
        weight_rom[2844] = 20;
        weight_rom[2845] = 27;
        weight_rom[2846] = 14;
        weight_rom[2847] = 9;
        weight_rom[2848] = 3;
        weight_rom[2849] = 20;
        weight_rom[2850] = -2;
        weight_rom[2851] = 18;
        weight_rom[2852] = -10;
        weight_rom[2853] = -85;
        weight_rom[2854] = -80;
        weight_rom[2855] = 3;
        weight_rom[2856] = -2;
        weight_rom[2857] = 3;
        weight_rom[2858] = -6;
        weight_rom[2859] = 36;
        weight_rom[2860] = -2;
        weight_rom[2861] = -5;
        weight_rom[2862] = 17;
        weight_rom[2863] = 2;
        weight_rom[2864] = -7;
        weight_rom[2865] = -16;
        weight_rom[2866] = -29;
        weight_rom[2867] = -15;
        weight_rom[2868] = -23;
        weight_rom[2869] = -11;
        weight_rom[2870] = -8;
        weight_rom[2871] = 14;
        weight_rom[2872] = 22;
        weight_rom[2873] = 13;
        weight_rom[2874] = 11;
        weight_rom[2875] = 9;
        weight_rom[2876] = 8;
        weight_rom[2877] = 12;
        weight_rom[2878] = -5;
        weight_rom[2879] = -15;
        weight_rom[2880] = -44;
        weight_rom[2881] = -93;
        weight_rom[2882] = -23;
        weight_rom[2883] = -15;
        weight_rom[2884] = 0;
        weight_rom[2885] = 6;
        weight_rom[2886] = 3;
        weight_rom[2887] = 37;
        weight_rom[2888] = -12;
        weight_rom[2889] = 16;
        weight_rom[2890] = -1;
        weight_rom[2891] = 1;
        weight_rom[2892] = -2;
        weight_rom[2893] = -13;
        weight_rom[2894] = -24;
        weight_rom[2895] = -32;
        weight_rom[2896] = -35;
        weight_rom[2897] = -32;
        weight_rom[2898] = -11;
        weight_rom[2899] = 0;
        weight_rom[2900] = 2;
        weight_rom[2901] = 9;
        weight_rom[2902] = 13;
        weight_rom[2903] = 10;
        weight_rom[2904] = -9;
        weight_rom[2905] = 0;
        weight_rom[2906] = -17;
        weight_rom[2907] = -10;
        weight_rom[2908] = -18;
        weight_rom[2909] = -68;
        weight_rom[2910] = -42;
        weight_rom[2911] = 1;
        weight_rom[2912] = -3;
        weight_rom[2913] = -25;
        weight_rom[2914] = 3;
        weight_rom[2915] = 22;
        weight_rom[2916] = -7;
        weight_rom[2917] = -17;
        weight_rom[2918] = -1;
        weight_rom[2919] = -5;
        weight_rom[2920] = -11;
        weight_rom[2921] = -8;
        weight_rom[2922] = -28;
        weight_rom[2923] = -28;
        weight_rom[2924] = -37;
        weight_rom[2925] = -19;
        weight_rom[2926] = -3;
        weight_rom[2927] = 3;
        weight_rom[2928] = 6;
        weight_rom[2929] = 11;
        weight_rom[2930] = -6;
        weight_rom[2931] = 8;
        weight_rom[2932] = 8;
        weight_rom[2933] = -19;
        weight_rom[2934] = -19;
        weight_rom[2935] = -28;
        weight_rom[2936] = -29;
        weight_rom[2937] = -29;
        weight_rom[2938] = -37;
        weight_rom[2939] = 3;
        weight_rom[2940] = -1;
        weight_rom[2941] = 6;
        weight_rom[2942] = -5;
        weight_rom[2943] = -19;
        weight_rom[2944] = -20;
        weight_rom[2945] = -22;
        weight_rom[2946] = -11;
        weight_rom[2947] = -13;
        weight_rom[2948] = -6;
        weight_rom[2949] = -17;
        weight_rom[2950] = -14;
        weight_rom[2951] = -26;
        weight_rom[2952] = -15;
        weight_rom[2953] = -7;
        weight_rom[2954] = -7;
        weight_rom[2955] = -8;
        weight_rom[2956] = 4;
        weight_rom[2957] = -1;
        weight_rom[2958] = -2;
        weight_rom[2959] = 3;
        weight_rom[2960] = -4;
        weight_rom[2961] = -8;
        weight_rom[2962] = -11;
        weight_rom[2963] = -51;
        weight_rom[2964] = -15;
        weight_rom[2965] = -31;
        weight_rom[2966] = -22;
        weight_rom[2967] = -3;
        weight_rom[2968] = 3;
        weight_rom[2969] = 1;
        weight_rom[2970] = 1;
        weight_rom[2971] = -7;
        weight_rom[2972] = -10;
        weight_rom[2973] = -30;
        weight_rom[2974] = -36;
        weight_rom[2975] = -11;
        weight_rom[2976] = -19;
        weight_rom[2977] = -13;
        weight_rom[2978] = -9;
        weight_rom[2979] = 2;
        weight_rom[2980] = 4;
        weight_rom[2981] = -7;
        weight_rom[2982] = -1;
        weight_rom[2983] = 2;
        weight_rom[2984] = -1;
        weight_rom[2985] = 4;
        weight_rom[2986] = -7;
        weight_rom[2987] = 1;
        weight_rom[2988] = -16;
        weight_rom[2989] = -7;
        weight_rom[2990] = -7;
        weight_rom[2991] = 3;
        weight_rom[2992] = 2;
        weight_rom[2993] = -7;
        weight_rom[2994] = -14;
        weight_rom[2995] = 1;
        weight_rom[2996] = 1;
        weight_rom[2997] = 1;
        weight_rom[2998] = 35;
        weight_rom[2999] = 30;
        weight_rom[3000] = 30;
        weight_rom[3001] = -14;
        weight_rom[3002] = -6;
        weight_rom[3003] = 0;
        weight_rom[3004] = -3;
        weight_rom[3005] = -5;
        weight_rom[3006] = 2;
        weight_rom[3007] = 5;
        weight_rom[3008] = -5;
        weight_rom[3009] = -2;
        weight_rom[3010] = 0;
        weight_rom[3011] = -10;
        weight_rom[3012] = -13;
        weight_rom[3013] = -3;
        weight_rom[3014] = 9;
        weight_rom[3015] = 3;
        weight_rom[3016] = -9;
        weight_rom[3017] = -17;
        weight_rom[3018] = -18;
        weight_rom[3019] = -7;
        weight_rom[3020] = -2;
        weight_rom[3021] = -10;
        weight_rom[3022] = -6;
        weight_rom[3023] = 0;
        weight_rom[3024] = -1;
        weight_rom[3025] = -1;
        weight_rom[3026] = 8;
        weight_rom[3027] = 61;
        weight_rom[3028] = 46;
        weight_rom[3029] = 42;
        weight_rom[3030] = 31;
        weight_rom[3031] = 58;
        weight_rom[3032] = 28;
        weight_rom[3033] = 5;
        weight_rom[3034] = 18;
        weight_rom[3035] = 37;
        weight_rom[3036] = -4;
        weight_rom[3037] = 16;
        weight_rom[3038] = 2;
        weight_rom[3039] = 1;
        weight_rom[3040] = 14;
        weight_rom[3041] = 5;
        weight_rom[3042] = 4;
        weight_rom[3043] = 14;
        weight_rom[3044] = 19;
        weight_rom[3045] = 12;
        weight_rom[3046] = 9;
        weight_rom[3047] = 44;
        weight_rom[3048] = -17;
        weight_rom[3049] = -40;
        weight_rom[3050] = 0;
        weight_rom[3051] = 1;
        weight_rom[3052] = 3;
        weight_rom[3053] = 0;
        weight_rom[3054] = 2;
        weight_rom[3055] = -3;
        weight_rom[3056] = 40;
        weight_rom[3057] = 112;
        weight_rom[3058] = 68;
        weight_rom[3059] = 83;
        weight_rom[3060] = 78;
        weight_rom[3061] = 91;
        weight_rom[3062] = 87;
        weight_rom[3063] = 67;
        weight_rom[3064] = 67;
        weight_rom[3065] = 62;
        weight_rom[3066] = 55;
        weight_rom[3067] = 38;
        weight_rom[3068] = 66;
        weight_rom[3069] = 67;
        weight_rom[3070] = 85;
        weight_rom[3071] = 97;
        weight_rom[3072] = 100;
        weight_rom[3073] = 91;
        weight_rom[3074] = 56;
        weight_rom[3075] = 66;
        weight_rom[3076] = 43;
        weight_rom[3077] = 1;
        weight_rom[3078] = -3;
        weight_rom[3079] = 2;
        weight_rom[3080] = -3;
        weight_rom[3081] = 1;
        weight_rom[3082] = -1;
        weight_rom[3083] = -1;
        weight_rom[3084] = 47;
        weight_rom[3085] = 48;
        weight_rom[3086] = 62;
        weight_rom[3087] = 73;
        weight_rom[3088] = 84;
        weight_rom[3089] = 82;
        weight_rom[3090] = 71;
        weight_rom[3091] = 72;
        weight_rom[3092] = 76;
        weight_rom[3093] = 121;
        weight_rom[3094] = 126;
        weight_rom[3095] = 72;
        weight_rom[3096] = 127;
        weight_rom[3097] = 111;
        weight_rom[3098] = 99;
        weight_rom[3099] = 105;
        weight_rom[3100] = 87;
        weight_rom[3101] = 84;
        weight_rom[3102] = 48;
        weight_rom[3103] = 29;
        weight_rom[3104] = -2;
        weight_rom[3105] = -1;
        weight_rom[3106] = 2;
        weight_rom[3107] = -1;
        weight_rom[3108] = -1;
        weight_rom[3109] = 0;
        weight_rom[3110] = -1;
        weight_rom[3111] = -3;
        weight_rom[3112] = 1;
        weight_rom[3113] = -7;
        weight_rom[3114] = -13;
        weight_rom[3115] = 20;
        weight_rom[3116] = 9;
        weight_rom[3117] = 13;
        weight_rom[3118] = 31;
        weight_rom[3119] = 6;
        weight_rom[3120] = 13;
        weight_rom[3121] = -12;
        weight_rom[3122] = 31;
        weight_rom[3123] = 22;
        weight_rom[3124] = 5;
        weight_rom[3125] = -18;
        weight_rom[3126] = 20;
        weight_rom[3127] = -8;
        weight_rom[3128] = 12;
        weight_rom[3129] = 21;
        weight_rom[3130] = 33;
        weight_rom[3131] = -3;
        weight_rom[3132] = 3;
        weight_rom[3133] = 0;
        weight_rom[3134] = 1;
        weight_rom[3135] = 1;
        weight_rom[3136] = 0;
        weight_rom[3137] = 3;
        weight_rom[3138] = 3;
        weight_rom[3139] = 3;
        weight_rom[3140] = -2;
        weight_rom[3141] = -2;
        weight_rom[3142] = 3;
        weight_rom[3143] = 1;
        weight_rom[3144] = 2;
        weight_rom[3145] = -3;
        weight_rom[3146] = -3;
        weight_rom[3147] = 2;
        weight_rom[3148] = 1;
        weight_rom[3149] = -15;
        weight_rom[3150] = -26;
        weight_rom[3151] = 3;
        weight_rom[3152] = -3;
        weight_rom[3153] = 2;
        weight_rom[3154] = -1;
        weight_rom[3155] = -3;
        weight_rom[3156] = -3;
        weight_rom[3157] = 0;
        weight_rom[3158] = -2;
        weight_rom[3159] = 1;
        weight_rom[3160] = 1;
        weight_rom[3161] = -2;
        weight_rom[3162] = 1;
        weight_rom[3163] = 2;
        weight_rom[3164] = 1;
        weight_rom[3165] = -2;
        weight_rom[3166] = -2;
        weight_rom[3167] = 0;
        weight_rom[3168] = 2;
        weight_rom[3169] = 2;
        weight_rom[3170] = 15;
        weight_rom[3171] = -1;
        weight_rom[3172] = 22;
        weight_rom[3173] = 27;
        weight_rom[3174] = 31;
        weight_rom[3175] = -12;
        weight_rom[3176] = -14;
        weight_rom[3177] = 43;
        weight_rom[3178] = -4;
        weight_rom[3179] = -18;
        weight_rom[3180] = -43;
        weight_rom[3181] = 1;
        weight_rom[3182] = 45;
        weight_rom[3183] = 35;
        weight_rom[3184] = 33;
        weight_rom[3185] = 8;
        weight_rom[3186] = -3;
        weight_rom[3187] = -1;
        weight_rom[3188] = 1;
        weight_rom[3189] = 0;
        weight_rom[3190] = -3;
        weight_rom[3191] = -1;
        weight_rom[3192] = -3;
        weight_rom[3193] = 1;
        weight_rom[3194] = 0;
        weight_rom[3195] = 0;
        weight_rom[3196] = 19;
        weight_rom[3197] = -2;
        weight_rom[3198] = 32;
        weight_rom[3199] = 28;
        weight_rom[3200] = 41;
        weight_rom[3201] = 22;
        weight_rom[3202] = 38;
        weight_rom[3203] = 31;
        weight_rom[3204] = 20;
        weight_rom[3205] = -3;
        weight_rom[3206] = 39;
        weight_rom[3207] = 39;
        weight_rom[3208] = 15;
        weight_rom[3209] = 5;
        weight_rom[3210] = 17;
        weight_rom[3211] = 22;
        weight_rom[3212] = 50;
        weight_rom[3213] = 15;
        weight_rom[3214] = 41;
        weight_rom[3215] = 55;
        weight_rom[3216] = 24;
        weight_rom[3217] = 10;
        weight_rom[3218] = 3;
        weight_rom[3219] = -3;
        weight_rom[3220] = -2;
        weight_rom[3221] = 3;
        weight_rom[3222] = 11;
        weight_rom[3223] = 1;
        weight_rom[3224] = -2;
        weight_rom[3225] = -23;
        weight_rom[3226] = 23;
        weight_rom[3227] = 27;
        weight_rom[3228] = -4;
        weight_rom[3229] = 31;
        weight_rom[3230] = 17;
        weight_rom[3231] = 0;
        weight_rom[3232] = -4;
        weight_rom[3233] = 6;
        weight_rom[3234] = -6;
        weight_rom[3235] = 4;
        weight_rom[3236] = 2;
        weight_rom[3237] = 14;
        weight_rom[3238] = 19;
        weight_rom[3239] = 20;
        weight_rom[3240] = 9;
        weight_rom[3241] = 36;
        weight_rom[3242] = 43;
        weight_rom[3243] = 27;
        weight_rom[3244] = 26;
        weight_rom[3245] = -29;
        weight_rom[3246] = 0;
        weight_rom[3247] = -3;
        weight_rom[3248] = 0;
        weight_rom[3249] = 1;
        weight_rom[3250] = -25;
        weight_rom[3251] = 2;
        weight_rom[3252] = 12;
        weight_rom[3253] = -10;
        weight_rom[3254] = 2;
        weight_rom[3255] = 7;
        weight_rom[3256] = 5;
        weight_rom[3257] = 11;
        weight_rom[3258] = 8;
        weight_rom[3259] = -1;
        weight_rom[3260] = 5;
        weight_rom[3261] = 7;
        weight_rom[3262] = 2;
        weight_rom[3263] = -8;
        weight_rom[3264] = 9;
        weight_rom[3265] = 12;
        weight_rom[3266] = -8;
        weight_rom[3267] = 15;
        weight_rom[3268] = 8;
        weight_rom[3269] = -4;
        weight_rom[3270] = 12;
        weight_rom[3271] = 12;
        weight_rom[3272] = -22;
        weight_rom[3273] = -17;
        weight_rom[3274] = -23;
        weight_rom[3275] = 1;
        weight_rom[3276] = -1;
        weight_rom[3277] = 2;
        weight_rom[3278] = -3;
        weight_rom[3279] = -28;
        weight_rom[3280] = -8;
        weight_rom[3281] = -26;
        weight_rom[3282] = -5;
        weight_rom[3283] = 2;
        weight_rom[3284] = 13;
        weight_rom[3285] = 13;
        weight_rom[3286] = 17;
        weight_rom[3287] = 8;
        weight_rom[3288] = 21;
        weight_rom[3289] = 13;
        weight_rom[3290] = 29;
        weight_rom[3291] = 14;
        weight_rom[3292] = 26;
        weight_rom[3293] = 26;
        weight_rom[3294] = 16;
        weight_rom[3295] = 21;
        weight_rom[3296] = 4;
        weight_rom[3297] = 2;
        weight_rom[3298] = -13;
        weight_rom[3299] = 7;
        weight_rom[3300] = -2;
        weight_rom[3301] = -5;
        weight_rom[3302] = 16;
        weight_rom[3303] = -2;
        weight_rom[3304] = -3;
        weight_rom[3305] = 0;
        weight_rom[3306] = -25;
        weight_rom[3307] = -44;
        weight_rom[3308] = -11;
        weight_rom[3309] = 10;
        weight_rom[3310] = -12;
        weight_rom[3311] = 24;
        weight_rom[3312] = 11;
        weight_rom[3313] = 14;
        weight_rom[3314] = -3;
        weight_rom[3315] = -5;
        weight_rom[3316] = -3;
        weight_rom[3317] = 4;
        weight_rom[3318] = 2;
        weight_rom[3319] = 9;
        weight_rom[3320] = -2;
        weight_rom[3321] = 1;
        weight_rom[3322] = -19;
        weight_rom[3323] = -6;
        weight_rom[3324] = -15;
        weight_rom[3325] = -19;
        weight_rom[3326] = -16;
        weight_rom[3327] = 26;
        weight_rom[3328] = 6;
        weight_rom[3329] = -6;
        weight_rom[3330] = -2;
        weight_rom[3331] = 14;
        weight_rom[3332] = 2;
        weight_rom[3333] = -27;
        weight_rom[3334] = 5;
        weight_rom[3335] = -42;
        weight_rom[3336] = 13;
        weight_rom[3337] = 2;
        weight_rom[3338] = 4;
        weight_rom[3339] = 2;
        weight_rom[3340] = 6;
        weight_rom[3341] = -1;
        weight_rom[3342] = -1;
        weight_rom[3343] = -6;
        weight_rom[3344] = -11;
        weight_rom[3345] = 2;
        weight_rom[3346] = 0;
        weight_rom[3347] = 13;
        weight_rom[3348] = 4;
        weight_rom[3349] = -15;
        weight_rom[3350] = -13;
        weight_rom[3351] = -19;
        weight_rom[3352] = -18;
        weight_rom[3353] = -10;
        weight_rom[3354] = 5;
        weight_rom[3355] = -3;
        weight_rom[3356] = 25;
        weight_rom[3357] = 7;
        weight_rom[3358] = 10;
        weight_rom[3359] = 6;
        weight_rom[3360] = -1;
        weight_rom[3361] = -36;
        weight_rom[3362] = -6;
        weight_rom[3363] = -19;
        weight_rom[3364] = -1;
        weight_rom[3365] = 12;
        weight_rom[3366] = -5;
        weight_rom[3367] = 0;
        weight_rom[3368] = 0;
        weight_rom[3369] = 4;
        weight_rom[3370] = -7;
        weight_rom[3371] = -7;
        weight_rom[3372] = -8;
        weight_rom[3373] = -14;
        weight_rom[3374] = -18;
        weight_rom[3375] = -8;
        weight_rom[3376] = -21;
        weight_rom[3377] = -21;
        weight_rom[3378] = -25;
        weight_rom[3379] = -12;
        weight_rom[3380] = -20;
        weight_rom[3381] = 0;
        weight_rom[3382] = -13;
        weight_rom[3383] = -13;
        weight_rom[3384] = 3;
        weight_rom[3385] = 4;
        weight_rom[3386] = -27;
        weight_rom[3387] = -27;
        weight_rom[3388] = -20;
        weight_rom[3389] = -42;
        weight_rom[3390] = -20;
        weight_rom[3391] = -40;
        weight_rom[3392] = -15;
        weight_rom[3393] = 6;
        weight_rom[3394] = 7;
        weight_rom[3395] = 10;
        weight_rom[3396] = -7;
        weight_rom[3397] = -1;
        weight_rom[3398] = -6;
        weight_rom[3399] = -13;
        weight_rom[3400] = -14;
        weight_rom[3401] = -17;
        weight_rom[3402] = -37;
        weight_rom[3403] = -33;
        weight_rom[3404] = -24;
        weight_rom[3405] = -16;
        weight_rom[3406] = -1;
        weight_rom[3407] = 5;
        weight_rom[3408] = 2;
        weight_rom[3409] = 13;
        weight_rom[3410] = -14;
        weight_rom[3411] = 16;
        weight_rom[3412] = -26;
        weight_rom[3413] = -48;
        weight_rom[3414] = -19;
        weight_rom[3415] = -27;
        weight_rom[3416] = -23;
        weight_rom[3417] = -38;
        weight_rom[3418] = -39;
        weight_rom[3419] = -48;
        weight_rom[3420] = -8;
        weight_rom[3421] = 2;
        weight_rom[3422] = 1;
        weight_rom[3423] = 0;
        weight_rom[3424] = 7;
        weight_rom[3425] = 6;
        weight_rom[3426] = 4;
        weight_rom[3427] = -10;
        weight_rom[3428] = -18;
        weight_rom[3429] = -38;
        weight_rom[3430] = -72;
        weight_rom[3431] = -59;
        weight_rom[3432] = -46;
        weight_rom[3433] = -10;
        weight_rom[3434] = -4;
        weight_rom[3435] = 13;
        weight_rom[3436] = 2;
        weight_rom[3437] = -4;
        weight_rom[3438] = 2;
        weight_rom[3439] = -28;
        weight_rom[3440] = -30;
        weight_rom[3441] = -67;
        weight_rom[3442] = -86;
        weight_rom[3443] = -26;
        weight_rom[3444] = -8;
        weight_rom[3445] = -43;
        weight_rom[3446] = -60;
        weight_rom[3447] = -34;
        weight_rom[3448] = -23;
        weight_rom[3449] = 10;
        weight_rom[3450] = 7;
        weight_rom[3451] = -7;
        weight_rom[3452] = 2;
        weight_rom[3453] = 7;
        weight_rom[3454] = 7;
        weight_rom[3455] = -5;
        weight_rom[3456] = -5;
        weight_rom[3457] = -49;
        weight_rom[3458] = -68;
        weight_rom[3459] = -44;
        weight_rom[3460] = -5;
        weight_rom[3461] = -3;
        weight_rom[3462] = 4;
        weight_rom[3463] = 23;
        weight_rom[3464] = 19;
        weight_rom[3465] = 16;
        weight_rom[3466] = 1;
        weight_rom[3467] = 22;
        weight_rom[3468] = 13;
        weight_rom[3469] = -49;
        weight_rom[3470] = -56;
        weight_rom[3471] = 26;
        weight_rom[3472] = -10;
        weight_rom[3473] = -12;
        weight_rom[3474] = -45;
        weight_rom[3475] = -50;
        weight_rom[3476] = -22;
        weight_rom[3477] = -15;
        weight_rom[3478] = -2;
        weight_rom[3479] = 2;
        weight_rom[3480] = 3;
        weight_rom[3481] = 18;
        weight_rom[3482] = 15;
        weight_rom[3483] = 26;
        weight_rom[3484] = 23;
        weight_rom[3485] = 11;
        weight_rom[3486] = -33;
        weight_rom[3487] = -9;
        weight_rom[3488] = 17;
        weight_rom[3489] = 17;
        weight_rom[3490] = 16;
        weight_rom[3491] = 32;
        weight_rom[3492] = 23;
        weight_rom[3493] = 35;
        weight_rom[3494] = 54;
        weight_rom[3495] = 86;
        weight_rom[3496] = 58;
        weight_rom[3497] = -30;
        weight_rom[3498] = -81;
        weight_rom[3499] = 30;
        weight_rom[3500] = 2;
        weight_rom[3501] = 4;
        weight_rom[3502] = -58;
        weight_rom[3503] = -35;
        weight_rom[3504] = -28;
        weight_rom[3505] = -5;
        weight_rom[3506] = 2;
        weight_rom[3507] = 8;
        weight_rom[3508] = 19;
        weight_rom[3509] = 24;
        weight_rom[3510] = 34;
        weight_rom[3511] = 34;
        weight_rom[3512] = 29;
        weight_rom[3513] = 25;
        weight_rom[3514] = 15;
        weight_rom[3515] = 26;
        weight_rom[3516] = 23;
        weight_rom[3517] = 26;
        weight_rom[3518] = 28;
        weight_rom[3519] = 22;
        weight_rom[3520] = 30;
        weight_rom[3521] = 28;
        weight_rom[3522] = 32;
        weight_rom[3523] = 54;
        weight_rom[3524] = 16;
        weight_rom[3525] = -19;
        weight_rom[3526] = -31;
        weight_rom[3527] = -8;
        weight_rom[3528] = -1;
        weight_rom[3529] = -20;
        weight_rom[3530] = 0;
        weight_rom[3531] = -13;
        weight_rom[3532] = 18;
        weight_rom[3533] = 20;
        weight_rom[3534] = 23;
        weight_rom[3535] = 31;
        weight_rom[3536] = 23;
        weight_rom[3537] = 28;
        weight_rom[3538] = 26;
        weight_rom[3539] = 56;
        weight_rom[3540] = 47;
        weight_rom[3541] = 30;
        weight_rom[3542] = 11;
        weight_rom[3543] = 11;
        weight_rom[3544] = 31;
        weight_rom[3545] = 18;
        weight_rom[3546] = 13;
        weight_rom[3547] = 18;
        weight_rom[3548] = -3;
        weight_rom[3549] = -10;
        weight_rom[3550] = 10;
        weight_rom[3551] = -15;
        weight_rom[3552] = -2;
        weight_rom[3553] = -6;
        weight_rom[3554] = -32;
        weight_rom[3555] = -1;
        weight_rom[3556] = -3;
        weight_rom[3557] = -24;
        weight_rom[3558] = -16;
        weight_rom[3559] = 32;
        weight_rom[3560] = 4;
        weight_rom[3561] = 12;
        weight_rom[3562] = 23;
        weight_rom[3563] = 28;
        weight_rom[3564] = 38;
        weight_rom[3565] = 28;
        weight_rom[3566] = 21;
        weight_rom[3567] = 38;
        weight_rom[3568] = 50;
        weight_rom[3569] = 33;
        weight_rom[3570] = 23;
        weight_rom[3571] = 16;
        weight_rom[3572] = 34;
        weight_rom[3573] = 25;
        weight_rom[3574] = -4;
        weight_rom[3575] = 0;
        weight_rom[3576] = -24;
        weight_rom[3577] = -21;
        weight_rom[3578] = -15;
        weight_rom[3579] = -22;
        weight_rom[3580] = -30;
        weight_rom[3581] = 28;
        weight_rom[3582] = 5;
        weight_rom[3583] = 15;
        weight_rom[3584] = -2;
        weight_rom[3585] = 2;
        weight_rom[3586] = -46;
        weight_rom[3587] = -7;
        weight_rom[3588] = -33;
        weight_rom[3589] = 23;
        weight_rom[3590] = 36;
        weight_rom[3591] = 43;
        weight_rom[3592] = 44;
        weight_rom[3593] = 32;
        weight_rom[3594] = 41;
        weight_rom[3595] = 48;
        weight_rom[3596] = 54;
        weight_rom[3597] = 21;
        weight_rom[3598] = 24;
        weight_rom[3599] = 31;
        weight_rom[3600] = 23;
        weight_rom[3601] = 20;
        weight_rom[3602] = 4;
        weight_rom[3603] = -13;
        weight_rom[3604] = -8;
        weight_rom[3605] = -3;
        weight_rom[3606] = -12;
        weight_rom[3607] = -5;
        weight_rom[3608] = 11;
        weight_rom[3609] = 42;
        weight_rom[3610] = -23;
        weight_rom[3611] = 2;
        weight_rom[3612] = -1;
        weight_rom[3613] = -4;
        weight_rom[3614] = 36;
        weight_rom[3615] = -25;
        weight_rom[3616] = -39;
        weight_rom[3617] = -5;
        weight_rom[3618] = 3;
        weight_rom[3619] = 29;
        weight_rom[3620] = 44;
        weight_rom[3621] = 52;
        weight_rom[3622] = 53;
        weight_rom[3623] = 54;
        weight_rom[3624] = 49;
        weight_rom[3625] = 28;
        weight_rom[3626] = 10;
        weight_rom[3627] = 13;
        weight_rom[3628] = 25;
        weight_rom[3629] = 16;
        weight_rom[3630] = 9;
        weight_rom[3631] = 2;
        weight_rom[3632] = -3;
        weight_rom[3633] = -7;
        weight_rom[3634] = 7;
        weight_rom[3635] = -13;
        weight_rom[3636] = -1;
        weight_rom[3637] = 35;
        weight_rom[3638] = -9;
        weight_rom[3639] = 3;
        weight_rom[3640] = 0;
        weight_rom[3641] = -4;
        weight_rom[3642] = 2;
        weight_rom[3643] = -19;
        weight_rom[3644] = -26;
        weight_rom[3645] = -6;
        weight_rom[3646] = 0;
        weight_rom[3647] = 36;
        weight_rom[3648] = 31;
        weight_rom[3649] = 48;
        weight_rom[3650] = 50;
        weight_rom[3651] = 37;
        weight_rom[3652] = 53;
        weight_rom[3653] = 14;
        weight_rom[3654] = 12;
        weight_rom[3655] = 11;
        weight_rom[3656] = 17;
        weight_rom[3657] = 9;
        weight_rom[3658] = 7;
        weight_rom[3659] = 5;
        weight_rom[3660] = 13;
        weight_rom[3661] = -5;
        weight_rom[3662] = -13;
        weight_rom[3663] = 21;
        weight_rom[3664] = 22;
        weight_rom[3665] = 16;
        weight_rom[3666] = 22;
        weight_rom[3667] = -6;
        weight_rom[3668] = -2;
        weight_rom[3669] = 0;
        weight_rom[3670] = 12;
        weight_rom[3671] = -45;
        weight_rom[3672] = -20;
        weight_rom[3673] = -16;
        weight_rom[3674] = 10;
        weight_rom[3675] = 17;
        weight_rom[3676] = 3;
        weight_rom[3677] = 10;
        weight_rom[3678] = 32;
        weight_rom[3679] = 32;
        weight_rom[3680] = 3;
        weight_rom[3681] = 3;
        weight_rom[3682] = 3;
        weight_rom[3683] = 16;
        weight_rom[3684] = 17;
        weight_rom[3685] = 14;
        weight_rom[3686] = 12;
        weight_rom[3687] = 13;
        weight_rom[3688] = 2;
        weight_rom[3689] = 15;
        weight_rom[3690] = 10;
        weight_rom[3691] = 16;
        weight_rom[3692] = -11;
        weight_rom[3693] = -20;
        weight_rom[3694] = 11;
        weight_rom[3695] = -22;
        weight_rom[3696] = 0;
        weight_rom[3697] = -26;
        weight_rom[3698] = 20;
        weight_rom[3699] = -22;
        weight_rom[3700] = -17;
        weight_rom[3701] = -20;
        weight_rom[3702] = -19;
        weight_rom[3703] = 15;
        weight_rom[3704] = -10;
        weight_rom[3705] = 5;
        weight_rom[3706] = 7;
        weight_rom[3707] = 5;
        weight_rom[3708] = 10;
        weight_rom[3709] = 5;
        weight_rom[3710] = 5;
        weight_rom[3711] = 30;
        weight_rom[3712] = 21;
        weight_rom[3713] = 10;
        weight_rom[3714] = 22;
        weight_rom[3715] = 6;
        weight_rom[3716] = 17;
        weight_rom[3717] = 18;
        weight_rom[3718] = 10;
        weight_rom[3719] = -3;
        weight_rom[3720] = -6;
        weight_rom[3721] = -8;
        weight_rom[3722] = 8;
        weight_rom[3723] = 1;
        weight_rom[3724] = -1;
        weight_rom[3725] = 14;
        weight_rom[3726] = 1;
        weight_rom[3727] = -34;
        weight_rom[3728] = -36;
        weight_rom[3729] = -26;
        weight_rom[3730] = -29;
        weight_rom[3731] = -10;
        weight_rom[3732] = -14;
        weight_rom[3733] = 6;
        weight_rom[3734] = 0;
        weight_rom[3735] = 5;
        weight_rom[3736] = 20;
        weight_rom[3737] = 17;
        weight_rom[3738] = 23;
        weight_rom[3739] = 6;
        weight_rom[3740] = 9;
        weight_rom[3741] = 24;
        weight_rom[3742] = 15;
        weight_rom[3743] = 17;
        weight_rom[3744] = 19;
        weight_rom[3745] = 16;
        weight_rom[3746] = 18;
        weight_rom[3747] = 31;
        weight_rom[3748] = 2;
        weight_rom[3749] = -19;
        weight_rom[3750] = 5;
        weight_rom[3751] = -1;
        weight_rom[3752] = -1;
        weight_rom[3753] = 0;
        weight_rom[3754] = 0;
        weight_rom[3755] = -3;
        weight_rom[3756] = -18;
        weight_rom[3757] = -44;
        weight_rom[3758] = -27;
        weight_rom[3759] = -19;
        weight_rom[3760] = -11;
        weight_rom[3761] = -16;
        weight_rom[3762] = 5;
        weight_rom[3763] = 5;
        weight_rom[3764] = 20;
        weight_rom[3765] = 24;
        weight_rom[3766] = 5;
        weight_rom[3767] = 2;
        weight_rom[3768] = -13;
        weight_rom[3769] = -7;
        weight_rom[3770] = 8;
        weight_rom[3771] = 9;
        weight_rom[3772] = 17;
        weight_rom[3773] = 31;
        weight_rom[3774] = 4;
        weight_rom[3775] = 9;
        weight_rom[3776] = 5;
        weight_rom[3777] = -16;
        weight_rom[3778] = -17;
        weight_rom[3779] = 2;
        weight_rom[3780] = -3;
        weight_rom[3781] = 3;
        weight_rom[3782] = -29;
        weight_rom[3783] = -13;
        weight_rom[3784] = -33;
        weight_rom[3785] = -33;
        weight_rom[3786] = -39;
        weight_rom[3787] = -35;
        weight_rom[3788] = 0;
        weight_rom[3789] = -9;
        weight_rom[3790] = -29;
        weight_rom[3791] = -8;
        weight_rom[3792] = -3;
        weight_rom[3793] = 11;
        weight_rom[3794] = 5;
        weight_rom[3795] = 0;
        weight_rom[3796] = 6;
        weight_rom[3797] = 4;
        weight_rom[3798] = 16;
        weight_rom[3799] = 30;
        weight_rom[3800] = 38;
        weight_rom[3801] = 53;
        weight_rom[3802] = 36;
        weight_rom[3803] = 48;
        weight_rom[3804] = -6;
        weight_rom[3805] = 12;
        weight_rom[3806] = -27;
        weight_rom[3807] = 0;
        weight_rom[3808] = 3;
        weight_rom[3809] = -3;
        weight_rom[3810] = -7;
        weight_rom[3811] = -75;
        weight_rom[3812] = -49;
        weight_rom[3813] = -52;
        weight_rom[3814] = -30;
        weight_rom[3815] = -22;
        weight_rom[3816] = -6;
        weight_rom[3817] = 5;
        weight_rom[3818] = 4;
        weight_rom[3819] = -2;
        weight_rom[3820] = -1;
        weight_rom[3821] = -10;
        weight_rom[3822] = 2;
        weight_rom[3823] = 2;
        weight_rom[3824] = 22;
        weight_rom[3825] = -3;
        weight_rom[3826] = 31;
        weight_rom[3827] = 12;
        weight_rom[3828] = 19;
        weight_rom[3829] = 18;
        weight_rom[3830] = 28;
        weight_rom[3831] = 14;
        weight_rom[3832] = -4;
        weight_rom[3833] = 37;
        weight_rom[3834] = -3;
        weight_rom[3835] = -1;
        weight_rom[3836] = 0;
        weight_rom[3837] = 2;
        weight_rom[3838] = -2;
        weight_rom[3839] = -15;
        weight_rom[3840] = -54;
        weight_rom[3841] = -45;
        weight_rom[3842] = -18;
        weight_rom[3843] = -19;
        weight_rom[3844] = -66;
        weight_rom[3845] = -48;
        weight_rom[3846] = -18;
        weight_rom[3847] = -34;
        weight_rom[3848] = -53;
        weight_rom[3849] = -27;
        weight_rom[3850] = -21;
        weight_rom[3851] = -17;
        weight_rom[3852] = -20;
        weight_rom[3853] = -28;
        weight_rom[3854] = -39;
        weight_rom[3855] = -46;
        weight_rom[3856] = -8;
        weight_rom[3857] = -28;
        weight_rom[3858] = -27;
        weight_rom[3859] = -25;
        weight_rom[3860] = -51;
        weight_rom[3861] = -1;
        weight_rom[3862] = -3;
        weight_rom[3863] = -2;
        weight_rom[3864] = 1;
        weight_rom[3865] = -3;
        weight_rom[3866] = -1;
        weight_rom[3867] = -3;
        weight_rom[3868] = 28;
        weight_rom[3869] = 14;
        weight_rom[3870] = 15;
        weight_rom[3871] = -10;
        weight_rom[3872] = -11;
        weight_rom[3873] = -39;
        weight_rom[3874] = -39;
        weight_rom[3875] = -33;
        weight_rom[3876] = -19;
        weight_rom[3877] = -48;
        weight_rom[3878] = -27;
        weight_rom[3879] = -47;
        weight_rom[3880] = -48;
        weight_rom[3881] = -56;
        weight_rom[3882] = -32;
        weight_rom[3883] = -45;
        weight_rom[3884] = -18;
        weight_rom[3885] = -21;
        weight_rom[3886] = -38;
        weight_rom[3887] = 5;
        weight_rom[3888] = -3;
        weight_rom[3889] = -1;
        weight_rom[3890] = 0;
        weight_rom[3891] = -2;
        weight_rom[3892] = -3;
        weight_rom[3893] = 0;
        weight_rom[3894] = 1;
        weight_rom[3895] = -1;
        weight_rom[3896] = -3;
        weight_rom[3897] = -18;
        weight_rom[3898] = -30;
        weight_rom[3899] = 0;
        weight_rom[3900] = -26;
        weight_rom[3901] = -32;
        weight_rom[3902] = -50;
        weight_rom[3903] = -12;
        weight_rom[3904] = -30;
        weight_rom[3905] = -47;
        weight_rom[3906] = -42;
        weight_rom[3907] = -21;
        weight_rom[3908] = 2;
        weight_rom[3909] = -26;
        weight_rom[3910] = -37;
        weight_rom[3911] = -10;
        weight_rom[3912] = 1;
        weight_rom[3913] = -9;
        weight_rom[3914] = 0;
        weight_rom[3915] = -2;
        weight_rom[3916] = -3;
        weight_rom[3917] = 3;
        weight_rom[3918] = 3;
        weight_rom[3919] = 0;
        weight_rom[3920] = 3;
        weight_rom[3921] = 2;
        weight_rom[3922] = 3;
        weight_rom[3923] = 0;
        weight_rom[3924] = 2;
        weight_rom[3925] = -3;
        weight_rom[3926] = 1;
        weight_rom[3927] = -2;
        weight_rom[3928] = -2;
        weight_rom[3929] = -2;
        weight_rom[3930] = -1;
        weight_rom[3931] = -1;
        weight_rom[3932] = 3;
        weight_rom[3933] = -15;
        weight_rom[3934] = -13;
        weight_rom[3935] = 0;
        weight_rom[3936] = 1;
        weight_rom[3937] = 0;
        weight_rom[3938] = 3;
        weight_rom[3939] = 2;
        weight_rom[3940] = 1;
        weight_rom[3941] = -3;
        weight_rom[3942] = 1;
        weight_rom[3943] = -3;
        weight_rom[3944] = -3;
        weight_rom[3945] = -2;
        weight_rom[3946] = 0;
        weight_rom[3947] = -3;
        weight_rom[3948] = -2;
        weight_rom[3949] = 1;
        weight_rom[3950] = 0;
        weight_rom[3951] = 2;
        weight_rom[3952] = 0;
        weight_rom[3953] = -1;
        weight_rom[3954] = -22;
        weight_rom[3955] = -37;
        weight_rom[3956] = -32;
        weight_rom[3957] = -37;
        weight_rom[3958] = -34;
        weight_rom[3959] = 6;
        weight_rom[3960] = -19;
        weight_rom[3961] = -50;
        weight_rom[3962] = -2;
        weight_rom[3963] = -48;
        weight_rom[3964] = 4;
        weight_rom[3965] = -52;
        weight_rom[3966] = -47;
        weight_rom[3967] = -37;
        weight_rom[3968] = -30;
        weight_rom[3969] = -28;
        weight_rom[3970] = -36;
        weight_rom[3971] = -25;
        weight_rom[3972] = -2;
        weight_rom[3973] = -1;
        weight_rom[3974] = 3;
        weight_rom[3975] = -3;
        weight_rom[3976] = 2;
        weight_rom[3977] = 0;
        weight_rom[3978] = 1;
        weight_rom[3979] = -1;
        weight_rom[3980] = -15;
        weight_rom[3981] = 0;
        weight_rom[3982] = -41;
        weight_rom[3983] = -41;
        weight_rom[3984] = -71;
        weight_rom[3985] = -90;
        weight_rom[3986] = -93;
        weight_rom[3987] = -93;
        weight_rom[3988] = -85;
        weight_rom[3989] = -94;
        weight_rom[3990] = -113;
        weight_rom[3991] = -100;
        weight_rom[3992] = -92;
        weight_rom[3993] = -76;
        weight_rom[3994] = -44;
        weight_rom[3995] = -49;
        weight_rom[3996] = -91;
        weight_rom[3997] = -63;
        weight_rom[3998] = -64;
        weight_rom[3999] = -56;
        weight_rom[4000] = -47;
        weight_rom[4001] = -36;
        weight_rom[4002] = -2;
        weight_rom[4003] = 0;
        weight_rom[4004] = 3;
        weight_rom[4005] = -3;
        weight_rom[4006] = -24;
        weight_rom[4007] = -2;
        weight_rom[4008] = -2;
        weight_rom[4009] = -32;
        weight_rom[4010] = -56;
        weight_rom[4011] = -86;
        weight_rom[4012] = -43;
        weight_rom[4013] = -50;
        weight_rom[4014] = -53;
        weight_rom[4015] = -50;
        weight_rom[4016] = -39;
        weight_rom[4017] = -51;
        weight_rom[4018] = -32;
        weight_rom[4019] = -52;
        weight_rom[4020] = -39;
        weight_rom[4021] = -25;
        weight_rom[4022] = -35;
        weight_rom[4023] = -37;
        weight_rom[4024] = -27;
        weight_rom[4025] = -11;
        weight_rom[4026] = -13;
        weight_rom[4027] = -10;
        weight_rom[4028] = -17;
        weight_rom[4029] = 2;
        weight_rom[4030] = 3;
        weight_rom[4031] = 1;
        weight_rom[4032] = 0;
        weight_rom[4033] = 0;
        weight_rom[4034] = 1;
        weight_rom[4035] = 2;
        weight_rom[4036] = 20;
        weight_rom[4037] = -27;
        weight_rom[4038] = -46;
        weight_rom[4039] = -18;
        weight_rom[4040] = -25;
        weight_rom[4041] = -2;
        weight_rom[4042] = -7;
        weight_rom[4043] = 9;
        weight_rom[4044] = 17;
        weight_rom[4045] = 1;
        weight_rom[4046] = 9;
        weight_rom[4047] = 26;
        weight_rom[4048] = 7;
        weight_rom[4049] = 2;
        weight_rom[4050] = 2;
        weight_rom[4051] = -10;
        weight_rom[4052] = -15;
        weight_rom[4053] = 6;
        weight_rom[4054] = -16;
        weight_rom[4055] = -7;
        weight_rom[4056] = 46;
        weight_rom[4057] = 33;
        weight_rom[4058] = 24;
        weight_rom[4059] = -2;
        weight_rom[4060] = -2;
        weight_rom[4061] = 1;
        weight_rom[4062] = 3;
        weight_rom[4063] = -16;
        weight_rom[4064] = -49;
        weight_rom[4065] = -32;
        weight_rom[4066] = -13;
        weight_rom[4067] = -13;
        weight_rom[4068] = 17;
        weight_rom[4069] = 8;
        weight_rom[4070] = 17;
        weight_rom[4071] = 42;
        weight_rom[4072] = 21;
        weight_rom[4073] = 29;
        weight_rom[4074] = 9;
        weight_rom[4075] = 15;
        weight_rom[4076] = 11;
        weight_rom[4077] = 25;
        weight_rom[4078] = -2;
        weight_rom[4079] = -11;
        weight_rom[4080] = 0;
        weight_rom[4081] = -9;
        weight_rom[4082] = -18;
        weight_rom[4083] = -17;
        weight_rom[4084] = 8;
        weight_rom[4085] = 43;
        weight_rom[4086] = -15;
        weight_rom[4087] = 2;
        weight_rom[4088] = -1;
        weight_rom[4089] = 2;
        weight_rom[4090] = 16;
        weight_rom[4091] = -36;
        weight_rom[4092] = -16;
        weight_rom[4093] = -16;
        weight_rom[4094] = -5;
        weight_rom[4095] = -10;
        weight_rom[4096] = 16;
        weight_rom[4097] = 8;
        weight_rom[4098] = 22;
        weight_rom[4099] = 25;
        weight_rom[4100] = 35;
        weight_rom[4101] = 25;
        weight_rom[4102] = 38;
        weight_rom[4103] = 45;
        weight_rom[4104] = 31;
        weight_rom[4105] = 37;
        weight_rom[4106] = 15;
        weight_rom[4107] = 17;
        weight_rom[4108] = 8;
        weight_rom[4109] = 12;
        weight_rom[4110] = 9;
        weight_rom[4111] = -17;
        weight_rom[4112] = 26;
        weight_rom[4113] = 71;
        weight_rom[4114] = 13;
        weight_rom[4115] = -19;
        weight_rom[4116] = -1;
        weight_rom[4117] = -34;
        weight_rom[4118] = -14;
        weight_rom[4119] = -23;
        weight_rom[4120] = -46;
        weight_rom[4121] = -20;
        weight_rom[4122] = 6;
        weight_rom[4123] = 17;
        weight_rom[4124] = 14;
        weight_rom[4125] = 31;
        weight_rom[4126] = 12;
        weight_rom[4127] = 30;
        weight_rom[4128] = 29;
        weight_rom[4129] = 31;
        weight_rom[4130] = 33;
        weight_rom[4131] = 51;
        weight_rom[4132] = 48;
        weight_rom[4133] = 36;
        weight_rom[4134] = 32;
        weight_rom[4135] = 17;
        weight_rom[4136] = 15;
        weight_rom[4137] = 12;
        weight_rom[4138] = 2;
        weight_rom[4139] = 31;
        weight_rom[4140] = 47;
        weight_rom[4141] = 51;
        weight_rom[4142] = -3;
        weight_rom[4143] = 0;
        weight_rom[4144] = 7;
        weight_rom[4145] = -16;
        weight_rom[4146] = -33;
        weight_rom[4147] = -35;
        weight_rom[4148] = -64;
        weight_rom[4149] = -6;
        weight_rom[4150] = 17;
        weight_rom[4151] = 5;
        weight_rom[4152] = 32;
        weight_rom[4153] = 25;
        weight_rom[4154] = 18;
        weight_rom[4155] = 15;
        weight_rom[4156] = 24;
        weight_rom[4157] = 27;
        weight_rom[4158] = 28;
        weight_rom[4159] = 24;
        weight_rom[4160] = 39;
        weight_rom[4161] = 16;
        weight_rom[4162] = 29;
        weight_rom[4163] = 17;
        weight_rom[4164] = 22;
        weight_rom[4165] = 24;
        weight_rom[4166] = 16;
        weight_rom[4167] = 46;
        weight_rom[4168] = 114;
        weight_rom[4169] = 76;
        weight_rom[4170] = 37;
        weight_rom[4171] = 16;
        weight_rom[4172] = -8;
        weight_rom[4173] = -18;
        weight_rom[4174] = -41;
        weight_rom[4175] = -28;
        weight_rom[4176] = -40;
        weight_rom[4177] = 10;
        weight_rom[4178] = 32;
        weight_rom[4179] = -1;
        weight_rom[4180] = 18;
        weight_rom[4181] = 14;
        weight_rom[4182] = 25;
        weight_rom[4183] = 24;
        weight_rom[4184] = 26;
        weight_rom[4185] = 24;
        weight_rom[4186] = 2;
        weight_rom[4187] = -19;
        weight_rom[4188] = 8;
        weight_rom[4189] = 21;
        weight_rom[4190] = 26;
        weight_rom[4191] = 29;
        weight_rom[4192] = 33;
        weight_rom[4193] = 16;
        weight_rom[4194] = 22;
        weight_rom[4195] = 44;
        weight_rom[4196] = 116;
        weight_rom[4197] = 88;
        weight_rom[4198] = 29;
        weight_rom[4199] = 19;
        weight_rom[4200] = -7;
        weight_rom[4201] = -13;
        weight_rom[4202] = 10;
        weight_rom[4203] = -49;
        weight_rom[4204] = 14;
        weight_rom[4205] = 11;
        weight_rom[4206] = 27;
        weight_rom[4207] = 13;
        weight_rom[4208] = 18;
        weight_rom[4209] = 36;
        weight_rom[4210] = 30;
        weight_rom[4211] = 32;
        weight_rom[4212] = 25;
        weight_rom[4213] = 2;
        weight_rom[4214] = -11;
        weight_rom[4215] = -29;
        weight_rom[4216] = -10;
        weight_rom[4217] = 1;
        weight_rom[4218] = 26;
        weight_rom[4219] = 24;
        weight_rom[4220] = 35;
        weight_rom[4221] = 24;
        weight_rom[4222] = 32;
        weight_rom[4223] = 61;
        weight_rom[4224] = 85;
        weight_rom[4225] = 56;
        weight_rom[4226] = 51;
        weight_rom[4227] = 33;
        weight_rom[4228] = 0;
        weight_rom[4229] = -16;
        weight_rom[4230] = -61;
        weight_rom[4231] = -38;
        weight_rom[4232] = -8;
        weight_rom[4233] = 3;
        weight_rom[4234] = 33;
        weight_rom[4235] = 36;
        weight_rom[4236] = 27;
        weight_rom[4237] = 22;
        weight_rom[4238] = 24;
        weight_rom[4239] = 15;
        weight_rom[4240] = 1;
        weight_rom[4241] = 3;
        weight_rom[4242] = -3;
        weight_rom[4243] = -20;
        weight_rom[4244] = -17;
        weight_rom[4245] = 14;
        weight_rom[4246] = 21;
        weight_rom[4247] = 14;
        weight_rom[4248] = 25;
        weight_rom[4249] = 28;
        weight_rom[4250] = 31;
        weight_rom[4251] = 21;
        weight_rom[4252] = 42;
        weight_rom[4253] = 37;
        weight_rom[4254] = 70;
        weight_rom[4255] = -27;
        weight_rom[4256] = 9;
        weight_rom[4257] = -34;
        weight_rom[4258] = -47;
        weight_rom[4259] = -25;
        weight_rom[4260] = 18;
        weight_rom[4261] = 30;
        weight_rom[4262] = 42;
        weight_rom[4263] = 17;
        weight_rom[4264] = 18;
        weight_rom[4265] = 11;
        weight_rom[4266] = 3;
        weight_rom[4267] = 10;
        weight_rom[4268] = -10;
        weight_rom[4269] = -1;
        weight_rom[4270] = -15;
        weight_rom[4271] = -19;
        weight_rom[4272] = -26;
        weight_rom[4273] = 5;
        weight_rom[4274] = 12;
        weight_rom[4275] = 24;
        weight_rom[4276] = 32;
        weight_rom[4277] = 18;
        weight_rom[4278] = 30;
        weight_rom[4279] = -9;
        weight_rom[4280] = -14;
        weight_rom[4281] = -15;
        weight_rom[4282] = 37;
        weight_rom[4283] = -25;
        weight_rom[4284] = 3;
        weight_rom[4285] = -25;
        weight_rom[4286] = -50;
        weight_rom[4287] = 22;
        weight_rom[4288] = 29;
        weight_rom[4289] = 37;
        weight_rom[4290] = 9;
        weight_rom[4291] = 30;
        weight_rom[4292] = 10;
        weight_rom[4293] = 11;
        weight_rom[4294] = 21;
        weight_rom[4295] = 13;
        weight_rom[4296] = 1;
        weight_rom[4297] = -7;
        weight_rom[4298] = -20;
        weight_rom[4299] = -15;
        weight_rom[4300] = -15;
        weight_rom[4301] = -7;
        weight_rom[4302] = 17;
        weight_rom[4303] = 22;
        weight_rom[4304] = 21;
        weight_rom[4305] = 8;
        weight_rom[4306] = 14;
        weight_rom[4307] = -10;
        weight_rom[4308] = -31;
        weight_rom[4309] = -14;
        weight_rom[4310] = -23;
        weight_rom[4311] = -40;
        weight_rom[4312] = -3;
        weight_rom[4313] = -11;
        weight_rom[4314] = -28;
        weight_rom[4315] = 1;
        weight_rom[4316] = 48;
        weight_rom[4317] = 3;
        weight_rom[4318] = 13;
        weight_rom[4319] = 18;
        weight_rom[4320] = -1;
        weight_rom[4321] = 6;
        weight_rom[4322] = 27;
        weight_rom[4323] = 1;
        weight_rom[4324] = -9;
        weight_rom[4325] = 19;
        weight_rom[4326] = -6;
        weight_rom[4327] = -18;
        weight_rom[4328] = -28;
        weight_rom[4329] = 16;
        weight_rom[4330] = 8;
        weight_rom[4331] = -1;
        weight_rom[4332] = -1;
        weight_rom[4333] = -2;
        weight_rom[4334] = -14;
        weight_rom[4335] = -18;
        weight_rom[4336] = 2;
        weight_rom[4337] = -28;
        weight_rom[4338] = -59;
        weight_rom[4339] = 0;
        weight_rom[4340] = 3;
        weight_rom[4341] = 11;
        weight_rom[4342] = -38;
        weight_rom[4343] = -18;
        weight_rom[4344] = 17;
        weight_rom[4345] = -12;
        weight_rom[4346] = -11;
        weight_rom[4347] = 14;
        weight_rom[4348] = 11;
        weight_rom[4349] = 23;
        weight_rom[4350] = 22;
        weight_rom[4351] = -3;
        weight_rom[4352] = -14;
        weight_rom[4353] = -7;
        weight_rom[4354] = -33;
        weight_rom[4355] = -16;
        weight_rom[4356] = -16;
        weight_rom[4357] = 4;
        weight_rom[4358] = 20;
        weight_rom[4359] = -6;
        weight_rom[4360] = -7;
        weight_rom[4361] = -23;
        weight_rom[4362] = -21;
        weight_rom[4363] = -7;
        weight_rom[4364] = -15;
        weight_rom[4365] = -32;
        weight_rom[4366] = -49;
        weight_rom[4367] = -25;
        weight_rom[4368] = 2;
        weight_rom[4369] = 3;
        weight_rom[4370] = -38;
        weight_rom[4371] = -30;
        weight_rom[4372] = -3;
        weight_rom[4373] = -25;
        weight_rom[4374] = 2;
        weight_rom[4375] = 6;
        weight_rom[4376] = 30;
        weight_rom[4377] = -3;
        weight_rom[4378] = -3;
        weight_rom[4379] = -7;
        weight_rom[4380] = 3;
        weight_rom[4381] = -19;
        weight_rom[4382] = -34;
        weight_rom[4383] = -16;
        weight_rom[4384] = -5;
        weight_rom[4385] = 15;
        weight_rom[4386] = 1;
        weight_rom[4387] = -15;
        weight_rom[4388] = -16;
        weight_rom[4389] = -27;
        weight_rom[4390] = -12;
        weight_rom[4391] = -2;
        weight_rom[4392] = -40;
        weight_rom[4393] = -62;
        weight_rom[4394] = -62;
        weight_rom[4395] = -39;
        weight_rom[4396] = 1;
        weight_rom[4397] = 1;
        weight_rom[4398] = -58;
        weight_rom[4399] = -39;
        weight_rom[4400] = -10;
        weight_rom[4401] = 4;
        weight_rom[4402] = 5;
        weight_rom[4403] = 3;
        weight_rom[4404] = 13;
        weight_rom[4405] = 18;
        weight_rom[4406] = 13;
        weight_rom[4407] = 16;
        weight_rom[4408] = 2;
        weight_rom[4409] = -22;
        weight_rom[4410] = -30;
        weight_rom[4411] = -4;
        weight_rom[4412] = 12;
        weight_rom[4413] = 18;
        weight_rom[4414] = 12;
        weight_rom[4415] = -11;
        weight_rom[4416] = 1;
        weight_rom[4417] = -9;
        weight_rom[4418] = -1;
        weight_rom[4419] = -5;
        weight_rom[4420] = 25;
        weight_rom[4421] = -31;
        weight_rom[4422] = -50;
        weight_rom[4423] = 3;
        weight_rom[4424] = -1;
        weight_rom[4425] = -3;
        weight_rom[4426] = -52;
        weight_rom[4427] = -39;
        weight_rom[4428] = 4;
        weight_rom[4429] = 1;
        weight_rom[4430] = 22;
        weight_rom[4431] = 13;
        weight_rom[4432] = 23;
        weight_rom[4433] = 22;
        weight_rom[4434] = 26;
        weight_rom[4435] = 19;
        weight_rom[4436] = -15;
        weight_rom[4437] = -18;
        weight_rom[4438] = -30;
        weight_rom[4439] = -4;
        weight_rom[4440] = -2;
        weight_rom[4441] = -3;
        weight_rom[4442] = -2;
        weight_rom[4443] = 0;
        weight_rom[4444] = -3;
        weight_rom[4445] = -3;
        weight_rom[4446] = 10;
        weight_rom[4447] = -12;
        weight_rom[4448] = -21;
        weight_rom[4449] = -54;
        weight_rom[4450] = -52;
        weight_rom[4451] = -28;
        weight_rom[4452] = 0;
        weight_rom[4453] = -1;
        weight_rom[4454] = 23;
        weight_rom[4455] = -33;
        weight_rom[4456] = -7;
        weight_rom[4457] = 25;
        weight_rom[4458] = 30;
        weight_rom[4459] = 21;
        weight_rom[4460] = 24;
        weight_rom[4461] = 8;
        weight_rom[4462] = 15;
        weight_rom[4463] = -13;
        weight_rom[4464] = 0;
        weight_rom[4465] = -20;
        weight_rom[4466] = -17;
        weight_rom[4467] = -20;
        weight_rom[4468] = -24;
        weight_rom[4469] = -15;
        weight_rom[4470] = -12;
        weight_rom[4471] = -2;
        weight_rom[4472] = 3;
        weight_rom[4473] = -9;
        weight_rom[4474] = 17;
        weight_rom[4475] = 21;
        weight_rom[4476] = 9;
        weight_rom[4477] = -26;
        weight_rom[4478] = -53;
        weight_rom[4479] = -17;
        weight_rom[4480] = 2;
        weight_rom[4481] = 22;
        weight_rom[4482] = 10;
        weight_rom[4483] = -33;
        weight_rom[4484] = -22;
        weight_rom[4485] = 23;
        weight_rom[4486] = 21;
        weight_rom[4487] = 9;
        weight_rom[4488] = 17;
        weight_rom[4489] = -1;
        weight_rom[4490] = -5;
        weight_rom[4491] = -16;
        weight_rom[4492] = -10;
        weight_rom[4493] = -6;
        weight_rom[4494] = -23;
        weight_rom[4495] = -20;
        weight_rom[4496] = -15;
        weight_rom[4497] = -16;
        weight_rom[4498] = -21;
        weight_rom[4499] = -10;
        weight_rom[4500] = -12;
        weight_rom[4501] = 7;
        weight_rom[4502] = 33;
        weight_rom[4503] = 21;
        weight_rom[4504] = -17;
        weight_rom[4505] = -25;
        weight_rom[4506] = -34;
        weight_rom[4507] = 1;
        weight_rom[4508] = -1;
        weight_rom[4509] = -21;
        weight_rom[4510] = -43;
        weight_rom[4511] = -45;
        weight_rom[4512] = -4;
        weight_rom[4513] = 5;
        weight_rom[4514] = 18;
        weight_rom[4515] = 16;
        weight_rom[4516] = 2;
        weight_rom[4517] = 11;
        weight_rom[4518] = -9;
        weight_rom[4519] = 0;
        weight_rom[4520] = -1;
        weight_rom[4521] = -12;
        weight_rom[4522] = -11;
        weight_rom[4523] = -6;
        weight_rom[4524] = -13;
        weight_rom[4525] = -30;
        weight_rom[4526] = -16;
        weight_rom[4527] = -17;
        weight_rom[4528] = -7;
        weight_rom[4529] = 8;
        weight_rom[4530] = 23;
        weight_rom[4531] = -2;
        weight_rom[4532] = -18;
        weight_rom[4533] = -22;
        weight_rom[4534] = -14;
        weight_rom[4535] = 0;
        weight_rom[4536] = 2;
        weight_rom[4537] = -1;
        weight_rom[4538] = -43;
        weight_rom[4539] = -39;
        weight_rom[4540] = -21;
        weight_rom[4541] = -22;
        weight_rom[4542] = -6;
        weight_rom[4543] = 10;
        weight_rom[4544] = 14;
        weight_rom[4545] = 5;
        weight_rom[4546] = 5;
        weight_rom[4547] = 7;
        weight_rom[4548] = 15;
        weight_rom[4549] = 29;
        weight_rom[4550] = 12;
        weight_rom[4551] = 1;
        weight_rom[4552] = 14;
        weight_rom[4553] = -7;
        weight_rom[4554] = -6;
        weight_rom[4555] = -10;
        weight_rom[4556] = -13;
        weight_rom[4557] = 3;
        weight_rom[4558] = 19;
        weight_rom[4559] = 21;
        weight_rom[4560] = 10;
        weight_rom[4561] = 8;
        weight_rom[4562] = -22;
        weight_rom[4563] = 2;
        weight_rom[4564] = -3;
        weight_rom[4565] = 0;
        weight_rom[4566] = -35;
        weight_rom[4567] = 8;
        weight_rom[4568] = -22;
        weight_rom[4569] = -15;
        weight_rom[4570] = -27;
        weight_rom[4571] = -6;
        weight_rom[4572] = 1;
        weight_rom[4573] = 7;
        weight_rom[4574] = 30;
        weight_rom[4575] = 29;
        weight_rom[4576] = 37;
        weight_rom[4577] = 39;
        weight_rom[4578] = 36;
        weight_rom[4579] = 10;
        weight_rom[4580] = 17;
        weight_rom[4581] = 6;
        weight_rom[4582] = -14;
        weight_rom[4583] = -20;
        weight_rom[4584] = -21;
        weight_rom[4585] = 3;
        weight_rom[4586] = -2;
        weight_rom[4587] = 10;
        weight_rom[4588] = 14;
        weight_rom[4589] = 2;
        weight_rom[4590] = -24;
        weight_rom[4591] = -2;
        weight_rom[4592] = -2;
        weight_rom[4593] = -2;
        weight_rom[4594] = -22;
        weight_rom[4595] = 29;
        weight_rom[4596] = -12;
        weight_rom[4597] = 8;
        weight_rom[4598] = -18;
        weight_rom[4599] = -1;
        weight_rom[4600] = 14;
        weight_rom[4601] = 6;
        weight_rom[4602] = 18;
        weight_rom[4603] = 28;
        weight_rom[4604] = 31;
        weight_rom[4605] = 37;
        weight_rom[4606] = 17;
        weight_rom[4607] = 22;
        weight_rom[4608] = 13;
        weight_rom[4609] = 10;
        weight_rom[4610] = 11;
        weight_rom[4611] = 3;
        weight_rom[4612] = 9;
        weight_rom[4613] = -14;
        weight_rom[4614] = -6;
        weight_rom[4615] = 57;
        weight_rom[4616] = 1;
        weight_rom[4617] = -39;
        weight_rom[4618] = -1;
        weight_rom[4619] = -2;
        weight_rom[4620] = -3;
        weight_rom[4621] = -1;
        weight_rom[4622] = 2;
        weight_rom[4623] = 27;
        weight_rom[4624] = 23;
        weight_rom[4625] = 14;
        weight_rom[4626] = -19;
        weight_rom[4627] = 23;
        weight_rom[4628] = -6;
        weight_rom[4629] = 18;
        weight_rom[4630] = 20;
        weight_rom[4631] = 40;
        weight_rom[4632] = 25;
        weight_rom[4633] = 60;
        weight_rom[4634] = 27;
        weight_rom[4635] = 53;
        weight_rom[4636] = 81;
        weight_rom[4637] = 74;
        weight_rom[4638] = 72;
        weight_rom[4639] = 76;
        weight_rom[4640] = 80;
        weight_rom[4641] = 101;
        weight_rom[4642] = 36;
        weight_rom[4643] = 67;
        weight_rom[4644] = 44;
        weight_rom[4645] = 0;
        weight_rom[4646] = 2;
        weight_rom[4647] = -3;
        weight_rom[4648] = -2;
        weight_rom[4649] = 0;
        weight_rom[4650] = 1;
        weight_rom[4651] = -2;
        weight_rom[4652] = 50;
        weight_rom[4653] = 14;
        weight_rom[4654] = -13;
        weight_rom[4655] = -13;
        weight_rom[4656] = 17;
        weight_rom[4657] = 39;
        weight_rom[4658] = 54;
        weight_rom[4659] = 64;
        weight_rom[4660] = 77;
        weight_rom[4661] = 91;
        weight_rom[4662] = 104;
        weight_rom[4663] = 83;
        weight_rom[4664] = 87;
        weight_rom[4665] = 73;
        weight_rom[4666] = 63;
        weight_rom[4667] = 56;
        weight_rom[4668] = 84;
        weight_rom[4669] = 92;
        weight_rom[4670] = 41;
        weight_rom[4671] = 28;
        weight_rom[4672] = -3;
        weight_rom[4673] = -2;
        weight_rom[4674] = 1;
        weight_rom[4675] = -2;
        weight_rom[4676] = -2;
        weight_rom[4677] = 0;
        weight_rom[4678] = -3;
        weight_rom[4679] = 3;
        weight_rom[4680] = 3;
        weight_rom[4681] = -27;
        weight_rom[4682] = -40;
        weight_rom[4683] = 12;
        weight_rom[4684] = -8;
        weight_rom[4685] = -3;
        weight_rom[4686] = 23;
        weight_rom[4687] = 10;
        weight_rom[4688] = 7;
        weight_rom[4689] = -55;
        weight_rom[4690] = 12;
        weight_rom[4691] = -6;
        weight_rom[4692] = -17;
        weight_rom[4693] = -52;
        weight_rom[4694] = -5;
        weight_rom[4695] = -13;
        weight_rom[4696] = -1;
        weight_rom[4697] = 29;
        weight_rom[4698] = 1;
        weight_rom[4699] = 2;
        weight_rom[4700] = 3;
        weight_rom[4701] = -2;
        weight_rom[4702] = 1;
        weight_rom[4703] = -1;
        weight_rom[4704] = -89;
        weight_rom[4705] = 127;
        weight_rom[4706] = 31;
        weight_rom[4707] = 103;
        weight_rom[4708] = -28;
        weight_rom[4709] = 72;
        weight_rom[4710] = -66;
        weight_rom[4711] = 1;
        weight_rom[4712] = 55;
        weight_rom[4713] = -86;
        weight_rom[4714] = -15;
        weight_rom[4715] = 82;
        weight_rom[4716] = 111;
        weight_rom[4717] = -15;
        weight_rom[4718] = -68;
        weight_rom[4719] = -20;
        weight_rom[4720] = -27;
        weight_rom[4721] = -91;
        weight_rom[4722] = 31;
        weight_rom[4723] = 72;
        weight_rom[4724] = 25;
        weight_rom[4725] = -75;
        weight_rom[4726] = 22;
        weight_rom[4727] = -34;
        weight_rom[4728] = 27;
        weight_rom[4729] = -6;
        weight_rom[4730] = 55;
        weight_rom[4731] = 67;
        weight_rom[4732] = -59;
        weight_rom[4733] = -24;
        weight_rom[4734] = -110;
        weight_rom[4735] = -27;
        weight_rom[4736] = -72;
        weight_rom[4737] = 57;
        weight_rom[4738] = 72;
        weight_rom[4739] = 8;
        weight_rom[4740] = -14;
        weight_rom[4741] = -127;
        weight_rom[4742] = 49;
        weight_rom[4743] = 14;
        weight_rom[4744] = -31;
        weight_rom[4745] = 62;
        weight_rom[4746] = -58;
        weight_rom[4747] = -50;
        weight_rom[4748] = 35;
        weight_rom[4749] = -59;
        weight_rom[4750] = 89;
        weight_rom[4751] = -24;
        weight_rom[4752] = -57;
        weight_rom[4753] = 121;
        weight_rom[4754] = -105;
        weight_rom[4755] = 46;
        weight_rom[4756] = -76;
        weight_rom[4757] = 41;
        weight_rom[4758] = 51;
        weight_rom[4759] = -61;
        weight_rom[4760] = -29;
        weight_rom[4761] = 3;
        weight_rom[4762] = 21;
        weight_rom[4763] = 47;
        weight_rom[4764] = -23;
        weight_rom[4765] = 11;
        weight_rom[4766] = -95;
        weight_rom[4767] = 60;
        weight_rom[4768] = 6;
        weight_rom[4769] = 51;
        weight_rom[4770] = -44;
        weight_rom[4771] = 126;
        weight_rom[4772] = -65;
        weight_rom[4773] = -88;
        weight_rom[4774] = 23;
        weight_rom[4775] = 113;
        weight_rom[4776] = -1;
        weight_rom[4777] = 35;
        weight_rom[4778] = -125;
        weight_rom[4779] = -46;
    end

    // 主状态机和MAC单元
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            valid <= 0;
            digit_out <= 0;
            neuron_idx <= 0;
            input_idx <= 0;
            accumulator <= 0;
        end else begin
            case (state)
                IDLE: begin
                    valid <= 0;
                    digit_out <= 0;
                    neuron_idx <= 0;
                    input_idx <= 0;
                    if (start) begin
                        state <= LAYER1_COMPUTE;
                        // 初始化累加器为第一个神经元的偏置
                        accumulator <= $signed(weight_rom[4704]);
                    end
                end

                LAYER1_COMPUTE: begin
                    // MAC操作: accumulator += weight * input
                    // 读取Layer1权重: 地址 = neuron_idx * 784 + input_idx
                    accumulator <= accumulator + ($signed(weight_rom[neuron_idx * 784 + input_idx]) * $signed({31'b0, image_in[input_idx]}));

                    if (input_idx == 783) begin
                        // 当前神经元计算完成，进入激活
                        state <= LAYER1_ACTIVATE;
                        input_idx <= 0;
                    end else begin
                        // 继续计算下一个输入
                        input_idx <= input_idx + 1;
                    end
                end

                LAYER1_ACTIVATE: begin
                    // ReLU激活
                    if (accumulator < 0) begin
                        layer1_out[neuron_idx] <= 0;
                    end else begin
                        layer1_out[neuron_idx] <= accumulator;
                    end

                    if (neuron_idx == 5) begin
                        // Layer1完成，进入Layer2
                        state <= LAYER2_COMPUTE;
                        neuron_idx <= 0;
                        input_idx <= 0;
                        // 初始化为Layer2第一个神经元的偏置
                        accumulator <= $signed(weight_rom[4770]);
                    end else begin
                        // 计算下一个神经元
                        neuron_idx <= neuron_idx + 1;
                        input_idx <= 0;
                        state <= LAYER1_COMPUTE;
                        // 加载下一个神经元的偏置
                        accumulator <= $signed(weight_rom[4704 + neuron_idx + 1]);
                    end
                end

                LAYER2_COMPUTE: begin
                    // MAC操作: accumulator += (weight * layer1_out) >> 7
                    // 读取Layer2权重
                    accumulator <= accumulator + (($signed(weight_rom[4710 + neuron_idx * 6 + input_idx]) * layer1_out[input_idx]) >>> 7);

                    if (input_idx == 5) begin
                        // 当前神经元计算完成
                        layer2_out[neuron_idx] <= accumulator;

                        if (neuron_idx == 9) begin
                            // Layer2完成，进入argmax
                            state <= ARGMAX;
                        end else begin
                            // 计算下一个神经元
                            neuron_idx <= neuron_idx + 1;
                            input_idx <= 0;
                            // 加载下一个神经元的偏置
                            accumulator <= $signed(weight_rom[4770 + neuron_idx + 1]);
                        end
                    end else begin
                        // 继续计算下一个输入
                        input_idx <= input_idx + 1;
                    end
                end

                ARGMAX: begin
                    // 找到最大值的索引（使用串行比较减少组合逻辑）
                    if (layer2_out[0] >= layer2_out[1] && layer2_out[0] >= layer2_out[2] &&
                        layer2_out[0] >= layer2_out[3] && layer2_out[0] >= layer2_out[4] &&
                        layer2_out[0] >= layer2_out[5] && layer2_out[0] >= layer2_out[6] &&
                        layer2_out[0] >= layer2_out[7] && layer2_out[0] >= layer2_out[8] &&
                        layer2_out[0] >= layer2_out[9])
                        digit_out <= 0;
                    else if (layer2_out[1] >= layer2_out[2] && layer2_out[1] >= layer2_out[3] &&
                             layer2_out[1] >= layer2_out[4] && layer2_out[1] >= layer2_out[5] &&
                             layer2_out[1] >= layer2_out[6] && layer2_out[1] >= layer2_out[7] &&
                             layer2_out[1] >= layer2_out[8] && layer2_out[1] >= layer2_out[9])
                        digit_out <= 1;
                    else if (layer2_out[2] >= layer2_out[3] && layer2_out[2] >= layer2_out[4] &&
                             layer2_out[2] >= layer2_out[5] && layer2_out[2] >= layer2_out[6] &&
                             layer2_out[2] >= layer2_out[7] && layer2_out[2] >= layer2_out[8] &&
                             layer2_out[2] >= layer2_out[9])
                        digit_out <= 2;
                    else if (layer2_out[3] >= layer2_out[4] && layer2_out[3] >= layer2_out[5] &&
                             layer2_out[3] >= layer2_out[6] && layer2_out[3] >= layer2_out[7] &&
                             layer2_out[3] >= layer2_out[8] && layer2_out[3] >= layer2_out[9])
                        digit_out <= 3;
                    else if (layer2_out[4] >= layer2_out[5] && layer2_out[4] >= layer2_out[6] &&
                             layer2_out[4] >= layer2_out[7] && layer2_out[4] >= layer2_out[8] &&
                             layer2_out[4] >= layer2_out[9])
                        digit_out <= 4;
                    else if (layer2_out[5] >= layer2_out[6] && layer2_out[5] >= layer2_out[7] &&
                             layer2_out[5] >= layer2_out[8] && layer2_out[5] >= layer2_out[9])
                        digit_out <= 5;
                    else if (layer2_out[6] >= layer2_out[7] && layer2_out[6] >= layer2_out[8] &&
                             layer2_out[6] >= layer2_out[9])
                        digit_out <= 6;
                    else if (layer2_out[7] >= layer2_out[8] && layer2_out[7] >= layer2_out[9])
                        digit_out <= 7;
                    else if (layer2_out[8] >= layer2_out[9])
                        digit_out <= 8;
                    else
                        digit_out <= 9;

                    valid <= 1;
                    state <= DONE;
                end

                DONE: begin
                    // 保持结果直到下一次start
                    valid <= 1;
                    // 允许在DONE状态重新开始新的计算
                    if (start) begin
                        state <= LAYER1_COMPUTE;
                        neuron_idx <= 0;
                        input_idx <= 0;
                        valid <= 0;
                        digit_out <= 0;
                        // 初始化累加器为第一个神经元的偏置
                        accumulator <= $signed(weight_rom[4704]);
                    end
                end

                default: begin
                    state <= IDLE;
                end
            endcase
        end
    end

endmodule
