// MNIST手写数字识别模型 - Int8量化版本（串行计算架构）
// MNIST手写数字识别模型 - Int8量化版本（高度优化串行架构）
// 极致优化：3个隐藏神经元，24位累加器，最小化逻辑资源
// 网络结构: 784 → 3 → 10
// 输入: 28x28二值图像 (784位)
// 输出: 预测数字 (0-9)
// 时钟周期: ~2395 cycles
// ROM大小: 2395 bytes
// 优化目标: LUT < 6,272

module mnist_model(
    input wire clk,
    input wire rst,
    input wire [783:0] image_in,
    input wire start,
    output reg [3:0] digit_out,
    output reg valid
);

    // 紧凑状态机 (2位足够5个状态)
    localparam IDLE = 2'd0;
    localparam LAYER1 = 2'd1;
    localparam LAYER2 = 2'd2;
    localparam ARGMAX = 2'd3;

    reg [1:0] state;
    reg [3:0] neuron_idx;    // 神经元索引 (0-9)
    reg [9:0] input_idx;     // 输入索引 (0-783)
    reg layer1_done;         // Layer1计算完成标志

    // 24位累加器（减少寄存器使用）
    reg signed [23:0] accumulator;

    // 层输出存储（24位）
    reg signed [23:0] layer1_out [0:2];
    reg signed [23:0] layer2_out [0:9];

    // Argmax变量
    reg [3:0] max_idx;
    reg signed [23:0] max_val;

    // ROM: 权重和偏置 (2395字节)
    // 强制使用BRAM以节省LUT
    (* ram_style = "block" *)
    (* ramstyle = "M9K" *)
    (* syn_ramstyle = "block_ram" *)
    reg signed [7:0] weight_rom [0:2394];

    // 初始化ROM
    initial begin
        weight_rom[0] = 2;
        weight_rom[1] = 0;
        weight_rom[2] = 0;
        weight_rom[3] = 0;
        weight_rom[4] = -1;
        weight_rom[5] = -1;
        weight_rom[6] = 0;
        weight_rom[7] = -1;
        weight_rom[8] = 2;
        weight_rom[9] = 0;
        weight_rom[10] = -1;
        weight_rom[11] = -1;
        weight_rom[12] = -2;
        weight_rom[13] = -4;
        weight_rom[14] = 0;
        weight_rom[15] = 1;
        weight_rom[16] = -2;
        weight_rom[17] = 1;
        weight_rom[18] = 0;
        weight_rom[19] = 0;
        weight_rom[20] = 0;
        weight_rom[21] = 1;
        weight_rom[22] = -1;
        weight_rom[23] = 1;
        weight_rom[24] = 0;
        weight_rom[25] = 1;
        weight_rom[26] = 0;
        weight_rom[27] = 0;
        weight_rom[28] = 1;
        weight_rom[29] = -1;
        weight_rom[30] = -2;
        weight_rom[31] = -1;
        weight_rom[32] = 1;
        weight_rom[33] = 2;
        weight_rom[34] = -1;
        weight_rom[35] = -26;
        weight_rom[36] = -6;
        weight_rom[37] = -22;
        weight_rom[38] = -45;
        weight_rom[39] = -48;
        weight_rom[40] = -34;
        weight_rom[41] = -33;
        weight_rom[42] = 19;
        weight_rom[43] = 28;
        weight_rom[44] = -17;
        weight_rom[45] = -41;
        weight_rom[46] = -35;
        weight_rom[47] = -30;
        weight_rom[48] = -40;
        weight_rom[49] = -28;
        weight_rom[50] = -34;
        weight_rom[51] = -23;
        weight_rom[52] = 0;
        weight_rom[53] = -1;
        weight_rom[54] = 2;
        weight_rom[55] = 1;
        weight_rom[56] = 1;
        weight_rom[57] = 1;
        weight_rom[58] = 2;
        weight_rom[59] = -2;
        weight_rom[60] = -14;
        weight_rom[61] = -2;
        weight_rom[62] = -28;
        weight_rom[63] = -51;
        weight_rom[64] = -47;
        weight_rom[65] = -72;
        weight_rom[66] = -91;
        weight_rom[67] = -87;
        weight_rom[68] = -91;
        weight_rom[69] = -99;
        weight_rom[70] = -96;
        weight_rom[71] = -48;
        weight_rom[72] = -93;
        weight_rom[73] = -75;
        weight_rom[74] = -63;
        weight_rom[75] = -45;
        weight_rom[76] = -27;
        weight_rom[77] = -57;
        weight_rom[78] = -50;
        weight_rom[79] = -46;
        weight_rom[80] = -30;
        weight_rom[81] = -19;
        weight_rom[82] = -1;
        weight_rom[83] = 1;
        weight_rom[84] = 2;
        weight_rom[85] = 2;
        weight_rom[86] = 0;
        weight_rom[87] = 2;
        weight_rom[88] = -2;
        weight_rom[89] = 2;
        weight_rom[90] = -45;
        weight_rom[91] = -74;
        weight_rom[92] = -94;
        weight_rom[93] = -65;
        weight_rom[94] = -108;
        weight_rom[95] = -106;
        weight_rom[96] = -127;
        weight_rom[97] = -92;
        weight_rom[98] = -98;
        weight_rom[99] = -92;
        weight_rom[100] = -99;
        weight_rom[101] = -81;
        weight_rom[102] = -90;
        weight_rom[103] = -75;
        weight_rom[104] = -79;
        weight_rom[105] = -51;
        weight_rom[106] = -33;
        weight_rom[107] = -43;
        weight_rom[108] = -47;
        weight_rom[109] = -14;
        weight_rom[110] = -2;
        weight_rom[111] = -2;
        weight_rom[112] = 2;
        weight_rom[113] = 0;
        weight_rom[114] = 27;
        weight_rom[115] = 1;
        weight_rom[116] = -3;
        weight_rom[117] = -1;
        weight_rom[118] = -25;
        weight_rom[119] = -13;
        weight_rom[120] = -1;
        weight_rom[121] = -21;
        weight_rom[122] = -11;
        weight_rom[123] = -3;
        weight_rom[124] = 0;
        weight_rom[125] = -2;
        weight_rom[126] = -4;
        weight_rom[127] = -4;
        weight_rom[128] = -8;
        weight_rom[129] = -3;
        weight_rom[130] = -9;
        weight_rom[131] = 4;
        weight_rom[132] = 7;
        weight_rom[133] = 6;
        weight_rom[134] = 7;
        weight_rom[135] = 8;
        weight_rom[136] = -15;
        weight_rom[137] = -18;
        weight_rom[138] = 9;
        weight_rom[139] = 0;
        weight_rom[140] = -2;
        weight_rom[141] = -2;
        weight_rom[142] = 0;
        weight_rom[143] = 31;
        weight_rom[144] = -22;
        weight_rom[145] = -3;
        weight_rom[146] = -1;
        weight_rom[147] = -10;
        weight_rom[148] = 2;
        weight_rom[149] = -2;
        weight_rom[150] = -11;
        weight_rom[151] = -2;
        weight_rom[152] = 7;
        weight_rom[153] = 4;
        weight_rom[154] = 1;
        weight_rom[155] = -2;
        weight_rom[156] = -3;
        weight_rom[157] = -9;
        weight_rom[158] = -4;
        weight_rom[159] = 4;
        weight_rom[160] = -3;
        weight_rom[161] = -5;
        weight_rom[162] = 1;
        weight_rom[163] = 2;
        weight_rom[164] = -5;
        weight_rom[165] = -1;
        weight_rom[166] = -12;
        weight_rom[167] = 2;
        weight_rom[168] = -2;
        weight_rom[169] = -1;
        weight_rom[170] = -12;
        weight_rom[171] = -11;
        weight_rom[172] = 0;
        weight_rom[173] = 9;
        weight_rom[174] = 4;
        weight_rom[175] = 0;
        weight_rom[176] = -1;
        weight_rom[177] = 0;
        weight_rom[178] = -4;
        weight_rom[179] = 2;
        weight_rom[180] = -2;
        weight_rom[181] = 0;
        weight_rom[182] = 8;
        weight_rom[183] = 5;
        weight_rom[184] = 2;
        weight_rom[185] = 7;
        weight_rom[186] = 0;
        weight_rom[187] = -5;
        weight_rom[188] = 4;
        weight_rom[189] = -4;
        weight_rom[190] = -2;
        weight_rom[191] = 2;
        weight_rom[192] = -13;
        weight_rom[193] = -6;
        weight_rom[194] = 6;
        weight_rom[195] = -28;
        weight_rom[196] = -1;
        weight_rom[197] = -29;
        weight_rom[198] = 10;
        weight_rom[199] = 18;
        weight_rom[200] = 6;
        weight_rom[201] = -10;
        weight_rom[202] = 1;
        weight_rom[203] = 5;
        weight_rom[204] = -2;
        weight_rom[205] = 1;
        weight_rom[206] = 2;
        weight_rom[207] = -3;
        weight_rom[208] = 2;
        weight_rom[209] = 4;
        weight_rom[210] = 4;
        weight_rom[211] = 5;
        weight_rom[212] = 7;
        weight_rom[213] = 0;
        weight_rom[214] = 1;
        weight_rom[215] = -2;
        weight_rom[216] = 3;
        weight_rom[217] = -6;
        weight_rom[218] = -2;
        weight_rom[219] = -3;
        weight_rom[220] = 2;
        weight_rom[221] = -25;
        weight_rom[222] = -2;
        weight_rom[223] = 6;
        weight_rom[224] = 21;
        weight_rom[225] = -3;
        weight_rom[226] = 4;
        weight_rom[227] = 6;
        weight_rom[228] = 12;
        weight_rom[229] = -6;
        weight_rom[230] = -3;
        weight_rom[231] = 1;
        weight_rom[232] = 11;
        weight_rom[233] = -4;
        weight_rom[234] = -2;
        weight_rom[235] = -4;
        weight_rom[236] = 4;
        weight_rom[237] = 8;
        weight_rom[238] = 8;
        weight_rom[239] = 3;
        weight_rom[240] = -2;
        weight_rom[241] = -2;
        weight_rom[242] = 2;
        weight_rom[243] = -3;
        weight_rom[244] = -5;
        weight_rom[245] = 3;
        weight_rom[246] = -8;
        weight_rom[247] = -4;
        weight_rom[248] = -5;
        weight_rom[249] = -14;
        weight_rom[250] = 5;
        weight_rom[251] = 9;
        weight_rom[252] = 22;
        weight_rom[253] = 6;
        weight_rom[254] = 12;
        weight_rom[255] = 25;
        weight_rom[256] = 9;
        weight_rom[257] = 4;
        weight_rom[258] = 10;
        weight_rom[259] = 1;
        weight_rom[260] = -3;
        weight_rom[261] = 6;
        weight_rom[262] = 4;
        weight_rom[263] = 1;
        weight_rom[264] = 3;
        weight_rom[265] = 2;
        weight_rom[266] = 5;
        weight_rom[267] = 6;
        weight_rom[268] = 2;
        weight_rom[269] = 2;
        weight_rom[270] = -1;
        weight_rom[271] = 0;
        weight_rom[272] = 2;
        weight_rom[273] = -4;
        weight_rom[274] = -2;
        weight_rom[275] = -7;
        weight_rom[276] = -20;
        weight_rom[277] = -23;
        weight_rom[278] = 5;
        weight_rom[279] = 24;
        weight_rom[280] = 25;
        weight_rom[281] = 74;
        weight_rom[282] = 13;
        weight_rom[283] = 2;
        weight_rom[284] = -8;
        weight_rom[285] = -1;
        weight_rom[286] = 5;
        weight_rom[287] = 7;
        weight_rom[288] = 6;
        weight_rom[289] = 3;
        weight_rom[290] = 4;
        weight_rom[291] = 3;
        weight_rom[292] = 0;
        weight_rom[293] = -5;
        weight_rom[294] = 6;
        weight_rom[295] = 9;
        weight_rom[296] = 2;
        weight_rom[297] = -1;
        weight_rom[298] = 1;
        weight_rom[299] = 3;
        weight_rom[300] = -1;
        weight_rom[301] = 3;
        weight_rom[302] = 8;
        weight_rom[303] = -13;
        weight_rom[304] = -29;
        weight_rom[305] = -19;
        weight_rom[306] = -7;
        weight_rom[307] = -12;
        weight_rom[308] = 37;
        weight_rom[309] = 62;
        weight_rom[310] = 24;
        weight_rom[311] = -18;
        weight_rom[312] = -3;
        weight_rom[313] = 5;
        weight_rom[314] = 7;
        weight_rom[315] = 6;
        weight_rom[316] = 6;
        weight_rom[317] = 10;
        weight_rom[318] = 7;
        weight_rom[319] = 6;
        weight_rom[320] = -2;
        weight_rom[321] = -8;
        weight_rom[322] = 22;
        weight_rom[323] = 19;
        weight_rom[324] = 4;
        weight_rom[325] = 9;
        weight_rom[326] = 9;
        weight_rom[327] = 3;
        weight_rom[328] = 12;
        weight_rom[329] = 8;
        weight_rom[330] = 15;
        weight_rom[331] = -9;
        weight_rom[332] = -17;
        weight_rom[333] = -7;
        weight_rom[334] = -10;
        weight_rom[335] = 2;
        weight_rom[336] = 21;
        weight_rom[337] = 2;
        weight_rom[338] = 19;
        weight_rom[339] = -19;
        weight_rom[340] = 11;
        weight_rom[341] = -3;
        weight_rom[342] = 3;
        weight_rom[343] = 5;
        weight_rom[344] = 2;
        weight_rom[345] = 3;
        weight_rom[346] = -7;
        weight_rom[347] = -1;
        weight_rom[348] = -13;
        weight_rom[349] = -7;
        weight_rom[350] = 38;
        weight_rom[351] = 17;
        weight_rom[352] = 7;
        weight_rom[353] = 14;
        weight_rom[354] = 15;
        weight_rom[355] = 17;
        weight_rom[356] = 12;
        weight_rom[357] = 11;
        weight_rom[358] = 17;
        weight_rom[359] = 5;
        weight_rom[360] = -52;
        weight_rom[361] = -17;
        weight_rom[362] = -14;
        weight_rom[363] = 0;
        weight_rom[364] = 0;
        weight_rom[365] = -20;
        weight_rom[366] = 32;
        weight_rom[367] = -9;
        weight_rom[368] = 31;
        weight_rom[369] = 3;
        weight_rom[370] = 0;
        weight_rom[371] = 6;
        weight_rom[372] = 6;
        weight_rom[373] = 4;
        weight_rom[374] = -2;
        weight_rom[375] = -13;
        weight_rom[376] = -20;
        weight_rom[377] = 9;
        weight_rom[378] = 36;
        weight_rom[379] = 27;
        weight_rom[380] = 7;
        weight_rom[381] = 11;
        weight_rom[382] = 18;
        weight_rom[383] = 14;
        weight_rom[384] = 20;
        weight_rom[385] = 15;
        weight_rom[386] = -2;
        weight_rom[387] = -33;
        weight_rom[388] = -46;
        weight_rom[389] = -43;
        weight_rom[390] = -39;
        weight_rom[391] = 1;
        weight_rom[392] = 1;
        weight_rom[393] = 23;
        weight_rom[394] = -2;
        weight_rom[395] = 6;
        weight_rom[396] = 22;
        weight_rom[397] = -5;
        weight_rom[398] = 1;
        weight_rom[399] = -6;
        weight_rom[400] = -5;
        weight_rom[401] = -7;
        weight_rom[402] = -11;
        weight_rom[403] = -10;
        weight_rom[404] = -13;
        weight_rom[405] = 22;
        weight_rom[406] = 36;
        weight_rom[407] = 15;
        weight_rom[408] = 1;
        weight_rom[409] = 11;
        weight_rom[410] = 11;
        weight_rom[411] = 8;
        weight_rom[412] = -3;
        weight_rom[413] = -6;
        weight_rom[414] = -12;
        weight_rom[415] = -17;
        weight_rom[416] = -50;
        weight_rom[417] = -25;
        weight_rom[418] = -46;
        weight_rom[419] = 2;
        weight_rom[420] = 0;
        weight_rom[421] = 11;
        weight_rom[422] = -8;
        weight_rom[423] = 3;
        weight_rom[424] = 8;
        weight_rom[425] = -16;
        weight_rom[426] = 8;
        weight_rom[427] = -3;
        weight_rom[428] = -4;
        weight_rom[429] = -8;
        weight_rom[430] = -11;
        weight_rom[431] = -12;
        weight_rom[432] = -1;
        weight_rom[433] = 25;
        weight_rom[434] = 31;
        weight_rom[435] = 11;
        weight_rom[436] = 2;
        weight_rom[437] = 11;
        weight_rom[438] = 5;
        weight_rom[439] = -7;
        weight_rom[440] = -10;
        weight_rom[441] = -4;
        weight_rom[442] = -9;
        weight_rom[443] = -5;
        weight_rom[444] = -32;
        weight_rom[445] = -41;
        weight_rom[446] = -63;
        weight_rom[447] = -22;
        weight_rom[448] = 2;
        weight_rom[449] = -1;
        weight_rom[450] = -20;
        weight_rom[451] = 7;
        weight_rom[452] = 3;
        weight_rom[453] = -3;
        weight_rom[454] = 10;
        weight_rom[455] = 4;
        weight_rom[456] = 1;
        weight_rom[457] = -4;
        weight_rom[458] = 0;
        weight_rom[459] = 1;
        weight_rom[460] = 11;
        weight_rom[461] = 24;
        weight_rom[462] = 20;
        weight_rom[463] = 2;
        weight_rom[464] = 6;
        weight_rom[465] = 3;
        weight_rom[466] = -7;
        weight_rom[467] = -9;
        weight_rom[468] = -7;
        weight_rom[469] = -20;
        weight_rom[470] = -4;
        weight_rom[471] = -4;
        weight_rom[472] = -42;
        weight_rom[473] = -69;
        weight_rom[474] = -38;
        weight_rom[475] = 1;
        weight_rom[476] = 1;
        weight_rom[477] = 3;
        weight_rom[478] = -18;
        weight_rom[479] = -17;
        weight_rom[480] = -17;
        weight_rom[481] = -6;
        weight_rom[482] = -14;
        weight_rom[483] = 0;
        weight_rom[484] = 4;
        weight_rom[485] = 8;
        weight_rom[486] = 4;
        weight_rom[487] = 10;
        weight_rom[488] = 15;
        weight_rom[489] = 24;
        weight_rom[490] = 17;
        weight_rom[491] = 2;
        weight_rom[492] = 1;
        weight_rom[493] = -5;
        weight_rom[494] = -8;
        weight_rom[495] = -8;
        weight_rom[496] = -2;
        weight_rom[497] = 2;
        weight_rom[498] = -1;
        weight_rom[499] = -8;
        weight_rom[500] = -67;
        weight_rom[501] = -65;
        weight_rom[502] = -49;
        weight_rom[503] = 0;
        weight_rom[504] = 2;
        weight_rom[505] = 2;
        weight_rom[506] = -4;
        weight_rom[507] = -14;
        weight_rom[508] = -27;
        weight_rom[509] = -23;
        weight_rom[510] = -12;
        weight_rom[511] = -6;
        weight_rom[512] = -7;
        weight_rom[513] = 1;
        weight_rom[514] = 2;
        weight_rom[515] = 12;
        weight_rom[516] = 7;
        weight_rom[517] = 21;
        weight_rom[518] = 13;
        weight_rom[519] = -1;
        weight_rom[520] = -7;
        weight_rom[521] = -11;
        weight_rom[522] = -6;
        weight_rom[523] = -13;
        weight_rom[524] = 0;
        weight_rom[525] = -8;
        weight_rom[526] = -7;
        weight_rom[527] = -26;
        weight_rom[528] = -102;
        weight_rom[529] = -49;
        weight_rom[530] = 2;
        weight_rom[531] = 23;
        weight_rom[532] = -1;
        weight_rom[533] = 3;
        weight_rom[534] = 18;
        weight_rom[535] = -5;
        weight_rom[536] = -22;
        weight_rom[537] = -27;
        weight_rom[538] = -18;
        weight_rom[539] = -18;
        weight_rom[540] = -13;
        weight_rom[541] = -11;
        weight_rom[542] = -15;
        weight_rom[543] = -14;
        weight_rom[544] = -15;
        weight_rom[545] = -4;
        weight_rom[546] = -2;
        weight_rom[547] = -7;
        weight_rom[548] = -12;
        weight_rom[549] = -14;
        weight_rom[550] = -15;
        weight_rom[551] = -7;
        weight_rom[552] = -13;
        weight_rom[553] = -18;
        weight_rom[554] = -13;
        weight_rom[555] = -16;
        weight_rom[556] = -68;
        weight_rom[557] = -14;
        weight_rom[558] = -24;
        weight_rom[559] = -2;
        weight_rom[560] = 1;
        weight_rom[561] = -27;
        weight_rom[562] = 7;
        weight_rom[563] = -5;
        weight_rom[564] = -34;
        weight_rom[565] = -20;
        weight_rom[566] = -14;
        weight_rom[567] = -8;
        weight_rom[568] = -18;
        weight_rom[569] = -7;
        weight_rom[570] = -16;
        weight_rom[571] = -11;
        weight_rom[572] = -16;
        weight_rom[573] = -8;
        weight_rom[574] = -1;
        weight_rom[575] = -8;
        weight_rom[576] = -8;
        weight_rom[577] = -5;
        weight_rom[578] = -9;
        weight_rom[579] = -8;
        weight_rom[580] = -5;
        weight_rom[581] = -9;
        weight_rom[582] = -3;
        weight_rom[583] = -11;
        weight_rom[584] = -54;
        weight_rom[585] = 1;
        weight_rom[586] = -7;
        weight_rom[587] = -2;
        weight_rom[588] = -1;
        weight_rom[589] = 24;
        weight_rom[590] = 2;
        weight_rom[591] = -28;
        weight_rom[592] = -20;
        weight_rom[593] = -8;
        weight_rom[594] = 2;
        weight_rom[595] = -10;
        weight_rom[596] = -2;
        weight_rom[597] = -3;
        weight_rom[598] = 0;
        weight_rom[599] = -11;
        weight_rom[600] = -5;
        weight_rom[601] = -7;
        weight_rom[602] = -5;
        weight_rom[603] = -8;
        weight_rom[604] = -10;
        weight_rom[605] = -9;
        weight_rom[606] = -14;
        weight_rom[607] = -8;
        weight_rom[608] = -7;
        weight_rom[609] = -7;
        weight_rom[610] = -16;
        weight_rom[611] = -34;
        weight_rom[612] = -11;
        weight_rom[613] = 4;
        weight_rom[614] = -46;
        weight_rom[615] = 0;
        weight_rom[616] = 1;
        weight_rom[617] = -1;
        weight_rom[618] = -2;
        weight_rom[619] = -7;
        weight_rom[620] = -5;
        weight_rom[621] = 8;
        weight_rom[622] = -8;
        weight_rom[623] = 5;
        weight_rom[624] = 1;
        weight_rom[625] = -5;
        weight_rom[626] = -1;
        weight_rom[627] = -5;
        weight_rom[628] = -9;
        weight_rom[629] = -10;
        weight_rom[630] = -1;
        weight_rom[631] = 0;
        weight_rom[632] = -4;
        weight_rom[633] = 4;
        weight_rom[634] = -11;
        weight_rom[635] = -4;
        weight_rom[636] = -4;
        weight_rom[637] = -15;
        weight_rom[638] = -5;
        weight_rom[639] = 2;
        weight_rom[640] = 0;
        weight_rom[641] = 27;
        weight_rom[642] = 4;
        weight_rom[643] = -1;
        weight_rom[644] = -2;
        weight_rom[645] = -2;
        weight_rom[646] = -3;
        weight_rom[647] = -18;
        weight_rom[648] = -7;
        weight_rom[649] = -15;
        weight_rom[650] = -4;
        weight_rom[651] = -4;
        weight_rom[652] = 0;
        weight_rom[653] = -4;
        weight_rom[654] = -12;
        weight_rom[655] = -5;
        weight_rom[656] = -3;
        weight_rom[657] = 1;
        weight_rom[658] = 0;
        weight_rom[659] = -2;
        weight_rom[660] = 3;
        weight_rom[661] = 3;
        weight_rom[662] = 1;
        weight_rom[663] = -10;
        weight_rom[664] = -9;
        weight_rom[665] = -7;
        weight_rom[666] = -5;
        weight_rom[667] = 4;
        weight_rom[668] = -5;
        weight_rom[669] = -12;
        weight_rom[670] = 26;
        weight_rom[671] = 1;
        weight_rom[672] = 1;
        weight_rom[673] = -1;
        weight_rom[674] = -16;
        weight_rom[675] = -16;
        weight_rom[676] = -8;
        weight_rom[677] = 4;
        weight_rom[678] = -6;
        weight_rom[679] = -8;
        weight_rom[680] = -4;
        weight_rom[681] = -12;
        weight_rom[682] = -4;
        weight_rom[683] = -9;
        weight_rom[684] = -9;
        weight_rom[685] = -11;
        weight_rom[686] = -13;
        weight_rom[687] = -6;
        weight_rom[688] = -6;
        weight_rom[689] = -8;
        weight_rom[690] = 3;
        weight_rom[691] = 8;
        weight_rom[692] = 19;
        weight_rom[693] = 15;
        weight_rom[694] = -1;
        weight_rom[695] = 13;
        weight_rom[696] = -8;
        weight_rom[697] = -22;
        weight_rom[698] = 0;
        weight_rom[699] = -1;
        weight_rom[700] = 0;
        weight_rom[701] = 2;
        weight_rom[702] = 0;
        weight_rom[703] = -19;
        weight_rom[704] = -17;
        weight_rom[705] = 6;
        weight_rom[706] = -12;
        weight_rom[707] = 8;
        weight_rom[708] = -11;
        weight_rom[709] = 9;
        weight_rom[710] = -9;
        weight_rom[711] = 2;
        weight_rom[712] = -3;
        weight_rom[713] = 2;
        weight_rom[714] = 2;
        weight_rom[715] = -1;
        weight_rom[716] = 8;
        weight_rom[717] = 12;
        weight_rom[718] = 24;
        weight_rom[719] = 39;
        weight_rom[720] = 43;
        weight_rom[721] = 51;
        weight_rom[722] = -4;
        weight_rom[723] = 27;
        weight_rom[724] = 16;
        weight_rom[725] = -2;
        weight_rom[726] = 0;
        weight_rom[727] = 0;
        weight_rom[728] = 2;
        weight_rom[729] = 1;
        weight_rom[730] = 2;
        weight_rom[731] = 0;
        weight_rom[732] = 35;
        weight_rom[733] = 16;
        weight_rom[734] = 13;
        weight_rom[735] = 56;
        weight_rom[736] = 62;
        weight_rom[737] = 53;
        weight_rom[738] = 38;
        weight_rom[739] = 52;
        weight_rom[740] = 31;
        weight_rom[741] = 53;
        weight_rom[742] = 57;
        weight_rom[743] = 38;
        weight_rom[744] = 45;
        weight_rom[745] = 48;
        weight_rom[746] = 32;
        weight_rom[747] = 30;
        weight_rom[748] = 21;
        weight_rom[749] = 14;
        weight_rom[750] = 15;
        weight_rom[751] = 11;
        weight_rom[752] = -2;
        weight_rom[753] = 1;
        weight_rom[754] = 0;
        weight_rom[755] = 2;
        weight_rom[756] = 0;
        weight_rom[757] = -2;
        weight_rom[758] = -1;
        weight_rom[759] = -1;
        weight_rom[760] = -1;
        weight_rom[761] = 40;
        weight_rom[762] = 76;
        weight_rom[763] = 40;
        weight_rom[764] = 53;
        weight_rom[765] = 71;
        weight_rom[766] = 79;
        weight_rom[767] = 16;
        weight_rom[768] = 35;
        weight_rom[769] = 123;
        weight_rom[770] = 110;
        weight_rom[771] = 84;
        weight_rom[772] = 91;
        weight_rom[773] = 114;
        weight_rom[774] = 62;
        weight_rom[775] = 54;
        weight_rom[776] = 6;
        weight_rom[777] = 13;
        weight_rom[778] = 13;
        weight_rom[779] = 1;
        weight_rom[780] = 0;
        weight_rom[781] = -2;
        weight_rom[782] = 1;
        weight_rom[783] = 0;
        weight_rom[784] = 0;
        weight_rom[785] = -1;
        weight_rom[786] = -1;
        weight_rom[787] = 2;
        weight_rom[788] = 2;
        weight_rom[789] = 0;
        weight_rom[790] = 1;
        weight_rom[791] = -2;
        weight_rom[792] = 1;
        weight_rom[793] = 1;
        weight_rom[794] = -2;
        weight_rom[795] = 0;
        weight_rom[796] = 0;
        weight_rom[797] = -22;
        weight_rom[798] = -25;
        weight_rom[799] = 0;
        weight_rom[800] = 0;
        weight_rom[801] = 2;
        weight_rom[802] = -2;
        weight_rom[803] = -2;
        weight_rom[804] = 0;
        weight_rom[805] = 1;
        weight_rom[806] = 0;
        weight_rom[807] = -1;
        weight_rom[808] = -2;
        weight_rom[809] = 1;
        weight_rom[810] = 0;
        weight_rom[811] = -2;
        weight_rom[812] = 2;
        weight_rom[813] = -1;
        weight_rom[814] = 0;
        weight_rom[815] = 0;
        weight_rom[816] = 0;
        weight_rom[817] = 0;
        weight_rom[818] = 29;
        weight_rom[819] = 47;
        weight_rom[820] = 23;
        weight_rom[821] = 70;
        weight_rom[822] = 88;
        weight_rom[823] = 22;
        weight_rom[824] = 25;
        weight_rom[825] = 51;
        weight_rom[826] = -10;
        weight_rom[827] = 2;
        weight_rom[828] = -34;
        weight_rom[829] = 19;
        weight_rom[830] = 83;
        weight_rom[831] = 51;
        weight_rom[832] = 55;
        weight_rom[833] = 36;
        weight_rom[834] = 37;
        weight_rom[835] = 23;
        weight_rom[836] = 0;
        weight_rom[837] = -2;
        weight_rom[838] = 0;
        weight_rom[839] = -1;
        weight_rom[840] = 0;
        weight_rom[841] = -1;
        weight_rom[842] = 1;
        weight_rom[843] = 1;
        weight_rom[844] = 29;
        weight_rom[845] = -1;
        weight_rom[846] = 47;
        weight_rom[847] = 54;
        weight_rom[848] = 58;
        weight_rom[849] = 67;
        weight_rom[850] = 82;
        weight_rom[851] = 55;
        weight_rom[852] = 86;
        weight_rom[853] = 57;
        weight_rom[854] = 65;
        weight_rom[855] = 57;
        weight_rom[856] = 80;
        weight_rom[857] = 61;
        weight_rom[858] = 74;
        weight_rom[859] = 69;
        weight_rom[860] = 85;
        weight_rom[861] = 56;
        weight_rom[862] = 72;
        weight_rom[863] = 43;
        weight_rom[864] = 39;
        weight_rom[865] = -6;
        weight_rom[866] = 0;
        weight_rom[867] = 0;
        weight_rom[868] = 1;
        weight_rom[869] = -2;
        weight_rom[870] = 25;
        weight_rom[871] = -1;
        weight_rom[872] = -2;
        weight_rom[873] = -25;
        weight_rom[874] = 52;
        weight_rom[875] = 46;
        weight_rom[876] = 17;
        weight_rom[877] = 48;
        weight_rom[878] = 30;
        weight_rom[879] = 6;
        weight_rom[880] = 11;
        weight_rom[881] = 9;
        weight_rom[882] = 15;
        weight_rom[883] = 18;
        weight_rom[884] = 21;
        weight_rom[885] = 28;
        weight_rom[886] = 42;
        weight_rom[887] = 40;
        weight_rom[888] = 49;
        weight_rom[889] = 53;
        weight_rom[890] = 54;
        weight_rom[891] = 33;
        weight_rom[892] = 49;
        weight_rom[893] = -17;
        weight_rom[894] = 1;
        weight_rom[895] = 1;
        weight_rom[896] = 1;
        weight_rom[897] = 2;
        weight_rom[898] = -26;
        weight_rom[899] = -1;
        weight_rom[900] = 8;
        weight_rom[901] = -2;
        weight_rom[902] = 5;
        weight_rom[903] = 10;
        weight_rom[904] = 5;
        weight_rom[905] = -2;
        weight_rom[906] = -6;
        weight_rom[907] = -8;
        weight_rom[908] = -2;
        weight_rom[909] = -1;
        weight_rom[910] = 1;
        weight_rom[911] = -5;
        weight_rom[912] = -6;
        weight_rom[913] = -2;
        weight_rom[914] = -9;
        weight_rom[915] = -3;
        weight_rom[916] = -10;
        weight_rom[917] = -9;
        weight_rom[918] = 1;
        weight_rom[919] = 15;
        weight_rom[920] = 4;
        weight_rom[921] = -14;
        weight_rom[922] = -33;
        weight_rom[923] = -2;
        weight_rom[924] = -1;
        weight_rom[925] = 1;
        weight_rom[926] = 0;
        weight_rom[927] = -35;
        weight_rom[928] = -15;
        weight_rom[929] = -15;
        weight_rom[930] = -16;
        weight_rom[931] = -5;
        weight_rom[932] = -6;
        weight_rom[933] = -3;
        weight_rom[934] = -6;
        weight_rom[935] = -12;
        weight_rom[936] = -1;
        weight_rom[937] = -2;
        weight_rom[938] = 6;
        weight_rom[939] = 2;
        weight_rom[940] = 9;
        weight_rom[941] = 12;
        weight_rom[942] = 8;
        weight_rom[943] = 9;
        weight_rom[944] = 8;
        weight_rom[945] = -4;
        weight_rom[946] = -2;
        weight_rom[947] = 3;
        weight_rom[948] = -8;
        weight_rom[949] = 10;
        weight_rom[950] = 3;
        weight_rom[951] = 0;
        weight_rom[952] = -1;
        weight_rom[953] = 0;
        weight_rom[954] = -30;
        weight_rom[955] = -34;
        weight_rom[956] = -10;
        weight_rom[957] = 5;
        weight_rom[958] = -19;
        weight_rom[959] = -1;
        weight_rom[960] = -6;
        weight_rom[961] = -3;
        weight_rom[962] = -10;
        weight_rom[963] = -11;
        weight_rom[964] = -8;
        weight_rom[965] = -9;
        weight_rom[966] = -11;
        weight_rom[967] = -3;
        weight_rom[968] = -12;
        weight_rom[969] = -4;
        weight_rom[970] = -10;
        weight_rom[971] = -5;
        weight_rom[972] = -6;
        weight_rom[973] = -2;
        weight_rom[974] = 0;
        weight_rom[975] = 10;
        weight_rom[976] = 11;
        weight_rom[977] = -1;
        weight_rom[978] = -11;
        weight_rom[979] = 25;
        weight_rom[980] = -1;
        weight_rom[981] = -24;
        weight_rom[982] = -20;
        weight_rom[983] = -35;
        weight_rom[984] = -3;
        weight_rom[985] = -10;
        weight_rom[986] = -13;
        weight_rom[987] = -4;
        weight_rom[988] = 0;
        weight_rom[989] = -9;
        weight_rom[990] = -4;
        weight_rom[991] = -8;
        weight_rom[992] = -12;
        weight_rom[993] = -10;
        weight_rom[994] = -10;
        weight_rom[995] = -4;
        weight_rom[996] = -6;
        weight_rom[997] = -13;
        weight_rom[998] = -8;
        weight_rom[999] = -14;
        weight_rom[1000] = -5;
        weight_rom[1001] = -6;
        weight_rom[1002] = 4;
        weight_rom[1003] = 7;
        weight_rom[1004] = 17;
        weight_rom[1005] = -5;
        weight_rom[1006] = -13;
        weight_rom[1007] = 27;
        weight_rom[1008] = -3;
        weight_rom[1009] = -30;
        weight_rom[1010] = -14;
        weight_rom[1011] = -18;
        weight_rom[1012] = -10;
        weight_rom[1013] = -13;
        weight_rom[1014] = -6;
        weight_rom[1015] = -5;
        weight_rom[1016] = -1;
        weight_rom[1017] = 3;
        weight_rom[1018] = -3;
        weight_rom[1019] = -6;
        weight_rom[1020] = -9;
        weight_rom[1021] = -8;
        weight_rom[1022] = -11;
        weight_rom[1023] = -10;
        weight_rom[1024] = -14;
        weight_rom[1025] = -18;
        weight_rom[1026] = -10;
        weight_rom[1027] = -11;
        weight_rom[1028] = -10;
        weight_rom[1029] = 2;
        weight_rom[1030] = -4;
        weight_rom[1031] = -2;
        weight_rom[1032] = 20;
        weight_rom[1033] = -7;
        weight_rom[1034] = -11;
        weight_rom[1035] = 21;
        weight_rom[1036] = -20;
        weight_rom[1037] = -35;
        weight_rom[1038] = -37;
        weight_rom[1039] = -40;
        weight_rom[1040] = -7;
        weight_rom[1041] = -10;
        weight_rom[1042] = 0;
        weight_rom[1043] = 0;
        weight_rom[1044] = -1;
        weight_rom[1045] = 4;
        weight_rom[1046] = -2;
        weight_rom[1047] = -4;
        weight_rom[1048] = -8;
        weight_rom[1049] = -12;
        weight_rom[1050] = -21;
        weight_rom[1051] = -16;
        weight_rom[1052] = -18;
        weight_rom[1053] = -16;
        weight_rom[1054] = -9;
        weight_rom[1055] = -10;
        weight_rom[1056] = -6;
        weight_rom[1057] = -2;
        weight_rom[1058] = -3;
        weight_rom[1059] = 8;
        weight_rom[1060] = 13;
        weight_rom[1061] = -1;
        weight_rom[1062] = 8;
        weight_rom[1063] = -30;
        weight_rom[1064] = -17;
        weight_rom[1065] = -22;
        weight_rom[1066] = -33;
        weight_rom[1067] = -29;
        weight_rom[1068] = -3;
        weight_rom[1069] = -3;
        weight_rom[1070] = 2;
        weight_rom[1071] = 6;
        weight_rom[1072] = 6;
        weight_rom[1073] = 7;
        weight_rom[1074] = 9;
        weight_rom[1075] = 7;
        weight_rom[1076] = 4;
        weight_rom[1077] = -8;
        weight_rom[1078] = -21;
        weight_rom[1079] = -26;
        weight_rom[1080] = -29;
        weight_rom[1081] = -17;
        weight_rom[1082] = -15;
        weight_rom[1083] = -14;
        weight_rom[1084] = -15;
        weight_rom[1085] = -9;
        weight_rom[1086] = -7;
        weight_rom[1087] = -5;
        weight_rom[1088] = -6;
        weight_rom[1089] = 8;
        weight_rom[1090] = -14;
        weight_rom[1091] = -8;
        weight_rom[1092] = 1;
        weight_rom[1093] = -36;
        weight_rom[1094] = -49;
        weight_rom[1095] = -23;
        weight_rom[1096] = -9;
        weight_rom[1097] = 5;
        weight_rom[1098] = 1;
        weight_rom[1099] = 2;
        weight_rom[1100] = 7;
        weight_rom[1101] = 10;
        weight_rom[1102] = 10;
        weight_rom[1103] = 14;
        weight_rom[1104] = 14;
        weight_rom[1105] = 1;
        weight_rom[1106] = 0;
        weight_rom[1107] = -9;
        weight_rom[1108] = -6;
        weight_rom[1109] = -5;
        weight_rom[1110] = -5;
        weight_rom[1111] = -3;
        weight_rom[1112] = -4;
        weight_rom[1113] = 0;
        weight_rom[1114] = -9;
        weight_rom[1115] = -7;
        weight_rom[1116] = 8;
        weight_rom[1117] = 5;
        weight_rom[1118] = 18;
        weight_rom[1119] = 25;
        weight_rom[1120] = -5;
        weight_rom[1121] = -8;
        weight_rom[1122] = -22;
        weight_rom[1123] = -32;
        weight_rom[1124] = 2;
        weight_rom[1125] = -7;
        weight_rom[1126] = 3;
        weight_rom[1127] = 6;
        weight_rom[1128] = 3;
        weight_rom[1129] = 8;
        weight_rom[1130] = 5;
        weight_rom[1131] = 15;
        weight_rom[1132] = 10;
        weight_rom[1133] = 12;
        weight_rom[1134] = 13;
        weight_rom[1135] = 13;
        weight_rom[1136] = 3;
        weight_rom[1137] = 9;
        weight_rom[1138] = 9;
        weight_rom[1139] = 11;
        weight_rom[1140] = 2;
        weight_rom[1141] = 7;
        weight_rom[1142] = 3;
        weight_rom[1143] = 13;
        weight_rom[1144] = 14;
        weight_rom[1145] = -31;
        weight_rom[1146] = -69;
        weight_rom[1147] = 28;
        weight_rom[1148] = 1;
        weight_rom[1149] = 15;
        weight_rom[1150] = -44;
        weight_rom[1151] = -18;
        weight_rom[1152] = 0;
        weight_rom[1153] = -1;
        weight_rom[1154] = -4;
        weight_rom[1155] = 1;
        weight_rom[1156] = 5;
        weight_rom[1157] = 6;
        weight_rom[1158] = 4;
        weight_rom[1159] = 5;
        weight_rom[1160] = 6;
        weight_rom[1161] = 14;
        weight_rom[1162] = 32;
        weight_rom[1163] = 23;
        weight_rom[1164] = 3;
        weight_rom[1165] = 11;
        weight_rom[1166] = 16;
        weight_rom[1167] = 10;
        weight_rom[1168] = 9;
        weight_rom[1169] = 12;
        weight_rom[1170] = -8;
        weight_rom[1171] = -2;
        weight_rom[1172] = -10;
        weight_rom[1173] = -30;
        weight_rom[1174] = -33;
        weight_rom[1175] = -19;
        weight_rom[1176] = 0;
        weight_rom[1177] = -25;
        weight_rom[1178] = 10;
        weight_rom[1179] = 4;
        weight_rom[1180] = 28;
        weight_rom[1181] = 5;
        weight_rom[1182] = 7;
        weight_rom[1183] = 2;
        weight_rom[1184] = 4;
        weight_rom[1185] = 2;
        weight_rom[1186] = 0;
        weight_rom[1187] = 20;
        weight_rom[1188] = 11;
        weight_rom[1189] = 24;
        weight_rom[1190] = 35;
        weight_rom[1191] = 13;
        weight_rom[1192] = 8;
        weight_rom[1193] = 7;
        weight_rom[1194] = 3;
        weight_rom[1195] = 1;
        weight_rom[1196] = -4;
        weight_rom[1197] = -10;
        weight_rom[1198] = -6;
        weight_rom[1199] = -19;
        weight_rom[1200] = 4;
        weight_rom[1201] = -10;
        weight_rom[1202] = -15;
        weight_rom[1203] = 1;
        weight_rom[1204] = -1;
        weight_rom[1205] = -24;
        weight_rom[1206] = -6;
        weight_rom[1207] = 29;
        weight_rom[1208] = -9;
        weight_rom[1209] = -7;
        weight_rom[1210] = 7;
        weight_rom[1211] = 3;
        weight_rom[1212] = 4;
        weight_rom[1213] = -2;
        weight_rom[1214] = 3;
        weight_rom[1215] = 9;
        weight_rom[1216] = 14;
        weight_rom[1217] = 32;
        weight_rom[1218] = 35;
        weight_rom[1219] = 12;
        weight_rom[1220] = 8;
        weight_rom[1221] = 4;
        weight_rom[1222] = -6;
        weight_rom[1223] = -11;
        weight_rom[1224] = -19;
        weight_rom[1225] = -12;
        weight_rom[1226] = -7;
        weight_rom[1227] = -8;
        weight_rom[1228] = -16;
        weight_rom[1229] = 34;
        weight_rom[1230] = 15;
        weight_rom[1231] = -10;
        weight_rom[1232] = 0;
        weight_rom[1233] = 0;
        weight_rom[1234] = -34;
        weight_rom[1235] = -11;
        weight_rom[1236] = -20;
        weight_rom[1237] = 4;
        weight_rom[1238] = 15;
        weight_rom[1239] = 5;
        weight_rom[1240] = 5;
        weight_rom[1241] = 3;
        weight_rom[1242] = 12;
        weight_rom[1243] = 20;
        weight_rom[1244] = 28;
        weight_rom[1245] = 26;
        weight_rom[1246] = 32;
        weight_rom[1247] = 14;
        weight_rom[1248] = 7;
        weight_rom[1249] = -1;
        weight_rom[1250] = -15;
        weight_rom[1251] = -17;
        weight_rom[1252] = -8;
        weight_rom[1253] = -6;
        weight_rom[1254] = -6;
        weight_rom[1255] = -10;
        weight_rom[1256] = 9;
        weight_rom[1257] = 32;
        weight_rom[1258] = -12;
        weight_rom[1259] = -3;
        weight_rom[1260] = -1;
        weight_rom[1261] = 0;
        weight_rom[1262] = 30;
        weight_rom[1263] = -15;
        weight_rom[1264] = -14;
        weight_rom[1265] = -8;
        weight_rom[1266] = -5;
        weight_rom[1267] = 1;
        weight_rom[1268] = 4;
        weight_rom[1269] = 15;
        weight_rom[1270] = 20;
        weight_rom[1271] = 26;
        weight_rom[1272] = 26;
        weight_rom[1273] = 25;
        weight_rom[1274] = 24;
        weight_rom[1275] = 8;
        weight_rom[1276] = 2;
        weight_rom[1277] = -5;
        weight_rom[1278] = -7;
        weight_rom[1279] = -10;
        weight_rom[1280] = -3;
        weight_rom[1281] = -11;
        weight_rom[1282] = -6;
        weight_rom[1283] = -16;
        weight_rom[1284] = 4;
        weight_rom[1285] = 31;
        weight_rom[1286] = -4;
        weight_rom[1287] = 0;
        weight_rom[1288] = 0;
        weight_rom[1289] = 1;
        weight_rom[1290] = -27;
        weight_rom[1291] = 1;
        weight_rom[1292] = -15;
        weight_rom[1293] = -3;
        weight_rom[1294] = -7;
        weight_rom[1295] = 0;
        weight_rom[1296] = 6;
        weight_rom[1297] = 14;
        weight_rom[1298] = 25;
        weight_rom[1299] = 22;
        weight_rom[1300] = 26;
        weight_rom[1301] = 15;
        weight_rom[1302] = 16;
        weight_rom[1303] = 3;
        weight_rom[1304] = 5;
        weight_rom[1305] = -1;
        weight_rom[1306] = -2;
        weight_rom[1307] = -2;
        weight_rom[1308] = 4;
        weight_rom[1309] = -9;
        weight_rom[1310] = -5;
        weight_rom[1311] = 6;
        weight_rom[1312] = 17;
        weight_rom[1313] = 28;
        weight_rom[1314] = 25;
        weight_rom[1315] = -8;
        weight_rom[1316] = 1;
        weight_rom[1317] = 0;
        weight_rom[1318] = -24;
        weight_rom[1319] = -15;
        weight_rom[1320] = -11;
        weight_rom[1321] = -11;
        weight_rom[1322] = -3;
        weight_rom[1323] = -3;
        weight_rom[1324] = -2;
        weight_rom[1325] = 6;
        weight_rom[1326] = 18;
        weight_rom[1327] = 17;
        weight_rom[1328] = 3;
        weight_rom[1329] = 9;
        weight_rom[1330] = 11;
        weight_rom[1331] = 13;
        weight_rom[1332] = 8;
        weight_rom[1333] = 8;
        weight_rom[1334] = 6;
        weight_rom[1335] = 1;
        weight_rom[1336] = -3;
        weight_rom[1337] = 10;
        weight_rom[1338] = 2;
        weight_rom[1339] = 10;
        weight_rom[1340] = 19;
        weight_rom[1341] = 14;
        weight_rom[1342] = 13;
        weight_rom[1343] = 21;
        weight_rom[1344] = -1;
        weight_rom[1345] = -24;
        weight_rom[1346] = 8;
        weight_rom[1347] = -16;
        weight_rom[1348] = -9;
        weight_rom[1349] = -6;
        weight_rom[1350] = -3;
        weight_rom[1351] = 5;
        weight_rom[1352] = 5;
        weight_rom[1353] = 6;
        weight_rom[1354] = 6;
        weight_rom[1355] = 0;
        weight_rom[1356] = 0;
        weight_rom[1357] = 0;
        weight_rom[1358] = 5;
        weight_rom[1359] = 12;
        weight_rom[1360] = 10;
        weight_rom[1361] = 4;
        weight_rom[1362] = 7;
        weight_rom[1363] = 3;
        weight_rom[1364] = 2;
        weight_rom[1365] = 0;
        weight_rom[1366] = 5;
        weight_rom[1367] = 14;
        weight_rom[1368] = 21;
        weight_rom[1369] = -1;
        weight_rom[1370] = 4;
        weight_rom[1371] = 0;
        weight_rom[1372] = -1;
        weight_rom[1373] = 25;
        weight_rom[1374] = -18;
        weight_rom[1375] = -16;
        weight_rom[1376] = -16;
        weight_rom[1377] = 1;
        weight_rom[1378] = 1;
        weight_rom[1379] = 3;
        weight_rom[1380] = -3;
        weight_rom[1381] = 3;
        weight_rom[1382] = -6;
        weight_rom[1383] = -2;
        weight_rom[1384] = 3;
        weight_rom[1385] = 1;
        weight_rom[1386] = 6;
        weight_rom[1387] = 0;
        weight_rom[1388] = -2;
        weight_rom[1389] = 10;
        weight_rom[1390] = 2;
        weight_rom[1391] = 5;
        weight_rom[1392] = 6;
        weight_rom[1393] = 4;
        weight_rom[1394] = 11;
        weight_rom[1395] = 32;
        weight_rom[1396] = 17;
        weight_rom[1397] = -20;
        weight_rom[1398] = 14;
        weight_rom[1399] = 1;
        weight_rom[1400] = -2;
        weight_rom[1401] = -2;
        weight_rom[1402] = -41;
        weight_rom[1403] = -1;
        weight_rom[1404] = 10;
        weight_rom[1405] = 5;
        weight_rom[1406] = -1;
        weight_rom[1407] = 0;
        weight_rom[1408] = -5;
        weight_rom[1409] = -12;
        weight_rom[1410] = -3;
        weight_rom[1411] = -3;
        weight_rom[1412] = -3;
        weight_rom[1413] = -2;
        weight_rom[1414] = -1;
        weight_rom[1415] = -4;
        weight_rom[1416] = -3;
        weight_rom[1417] = 2;
        weight_rom[1418] = 4;
        weight_rom[1419] = 5;
        weight_rom[1420] = 9;
        weight_rom[1421] = 10;
        weight_rom[1422] = 7;
        weight_rom[1423] = 13;
        weight_rom[1424] = 10;
        weight_rom[1425] = -18;
        weight_rom[1426] = -36;
        weight_rom[1427] = -1;
        weight_rom[1428] = 1;
        weight_rom[1429] = -1;
        weight_rom[1430] = -25;
        weight_rom[1431] = 2;
        weight_rom[1432] = -3;
        weight_rom[1433] = -18;
        weight_rom[1434] = -1;
        weight_rom[1435] = -11;
        weight_rom[1436] = 6;
        weight_rom[1437] = 4;
        weight_rom[1438] = -9;
        weight_rom[1439] = 0;
        weight_rom[1440] = 1;
        weight_rom[1441] = 3;
        weight_rom[1442] = 4;
        weight_rom[1443] = 3;
        weight_rom[1444] = 6;
        weight_rom[1445] = 3;
        weight_rom[1446] = 6;
        weight_rom[1447] = 11;
        weight_rom[1448] = 23;
        weight_rom[1449] = 19;
        weight_rom[1450] = 3;
        weight_rom[1451] = 2;
        weight_rom[1452] = -4;
        weight_rom[1453] = 5;
        weight_rom[1454] = -26;
        weight_rom[1455] = 1;
        weight_rom[1456] = 1;
        weight_rom[1457] = -1;
        weight_rom[1458] = 0;
        weight_rom[1459] = -62;
        weight_rom[1460] = -36;
        weight_rom[1461] = -50;
        weight_rom[1462] = -25;
        weight_rom[1463] = -17;
        weight_rom[1464] = -6;
        weight_rom[1465] = -3;
        weight_rom[1466] = 2;
        weight_rom[1467] = 3;
        weight_rom[1468] = 5;
        weight_rom[1469] = 2;
        weight_rom[1470] = 6;
        weight_rom[1471] = 6;
        weight_rom[1472] = 12;
        weight_rom[1473] = 1;
        weight_rom[1474] = 20;
        weight_rom[1475] = 18;
        weight_rom[1476] = 19;
        weight_rom[1477] = 7;
        weight_rom[1478] = 8;
        weight_rom[1479] = 7;
        weight_rom[1480] = -6;
        weight_rom[1481] = 8;
        weight_rom[1482] = 0;
        weight_rom[1483] = 0;
        weight_rom[1484] = 1;
        weight_rom[1485] = 1;
        weight_rom[1486] = -1;
        weight_rom[1487] = -3;
        weight_rom[1488] = -39;
        weight_rom[1489] = -18;
        weight_rom[1490] = -19;
        weight_rom[1491] = -8;
        weight_rom[1492] = -21;
        weight_rom[1493] = -17;
        weight_rom[1494] = -15;
        weight_rom[1495] = -22;
        weight_rom[1496] = -25;
        weight_rom[1497] = -20;
        weight_rom[1498] = -12;
        weight_rom[1499] = -18;
        weight_rom[1500] = -7;
        weight_rom[1501] = 3;
        weight_rom[1502] = -1;
        weight_rom[1503] = -2;
        weight_rom[1504] = 24;
        weight_rom[1505] = 10;
        weight_rom[1506] = 2;
        weight_rom[1507] = -20;
        weight_rom[1508] = -38;
        weight_rom[1509] = 0;
        weight_rom[1510] = 0;
        weight_rom[1511] = 0;
        weight_rom[1512] = 1;
        weight_rom[1513] = -1;
        weight_rom[1514] = 0;
        weight_rom[1515] = 1;
        weight_rom[1516] = 7;
        weight_rom[1517] = 12;
        weight_rom[1518] = 12;
        weight_rom[1519] = -16;
        weight_rom[1520] = -10;
        weight_rom[1521] = -3;
        weight_rom[1522] = 0;
        weight_rom[1523] = 5;
        weight_rom[1524] = 18;
        weight_rom[1525] = 6;
        weight_rom[1526] = 12;
        weight_rom[1527] = 8;
        weight_rom[1528] = 8;
        weight_rom[1529] = 9;
        weight_rom[1530] = 23;
        weight_rom[1531] = 9;
        weight_rom[1532] = 23;
        weight_rom[1533] = 10;
        weight_rom[1534] = -5;
        weight_rom[1535] = 13;
        weight_rom[1536] = 1;
        weight_rom[1537] = 0;
        weight_rom[1538] = 0;
        weight_rom[1539] = 1;
        weight_rom[1540] = -2;
        weight_rom[1541] = -1;
        weight_rom[1542] = -1;
        weight_rom[1543] = -2;
        weight_rom[1544] = 1;
        weight_rom[1545] = -25;
        weight_rom[1546] = -34;
        weight_rom[1547] = 2;
        weight_rom[1548] = -27;
        weight_rom[1549] = -30;
        weight_rom[1550] = -30;
        weight_rom[1551] = -1;
        weight_rom[1552] = -17;
        weight_rom[1553] = -38;
        weight_rom[1554] = -13;
        weight_rom[1555] = 9;
        weight_rom[1556] = -1;
        weight_rom[1557] = -21;
        weight_rom[1558] = -20;
        weight_rom[1559] = -19;
        weight_rom[1560] = 18;
        weight_rom[1561] = -1;
        weight_rom[1562] = -2;
        weight_rom[1563] = -1;
        weight_rom[1564] = 0;
        weight_rom[1565] = 1;
        weight_rom[1566] = 0;
        weight_rom[1567] = 1;
        weight_rom[1568] = 0;
        weight_rom[1569] = -2;
        weight_rom[1570] = 1;
        weight_rom[1571] = -1;
        weight_rom[1572] = 2;
        weight_rom[1573] = -1;
        weight_rom[1574] = 1;
        weight_rom[1575] = -2;
        weight_rom[1576] = -1;
        weight_rom[1577] = 1;
        weight_rom[1578] = 0;
        weight_rom[1579] = 1;
        weight_rom[1580] = 0;
        weight_rom[1581] = 20;
        weight_rom[1582] = 24;
        weight_rom[1583] = -1;
        weight_rom[1584] = -1;
        weight_rom[1585] = -2;
        weight_rom[1586] = 2;
        weight_rom[1587] = -1;
        weight_rom[1588] = 0;
        weight_rom[1589] = -1;
        weight_rom[1590] = 0;
        weight_rom[1591] = 0;
        weight_rom[1592] = -1;
        weight_rom[1593] = -1;
        weight_rom[1594] = 1;
        weight_rom[1595] = -1;
        weight_rom[1596] = -1;
        weight_rom[1597] = 2;
        weight_rom[1598] = 1;
        weight_rom[1599] = -2;
        weight_rom[1600] = -2;
        weight_rom[1601] = 1;
        weight_rom[1602] = -11;
        weight_rom[1603] = 10;
        weight_rom[1604] = 23;
        weight_rom[1605] = 21;
        weight_rom[1606] = 26;
        weight_rom[1607] = -10;
        weight_rom[1608] = -26;
        weight_rom[1609] = -10;
        weight_rom[1610] = 16;
        weight_rom[1611] = 3;
        weight_rom[1612] = 67;
        weight_rom[1613] = 11;
        weight_rom[1614] = -8;
        weight_rom[1615] = 23;
        weight_rom[1616] = -3;
        weight_rom[1617] = 24;
        weight_rom[1618] = 29;
        weight_rom[1619] = 16;
        weight_rom[1620] = 2;
        weight_rom[1621] = 0;
        weight_rom[1622] = 2;
        weight_rom[1623] = 0;
        weight_rom[1624] = -2;
        weight_rom[1625] = 0;
        weight_rom[1626] = 0;
        weight_rom[1627] = 2;
        weight_rom[1628] = -22;
        weight_rom[1629] = 0;
        weight_rom[1630] = -6;
        weight_rom[1631] = 0;
        weight_rom[1632] = 17;
        weight_rom[1633] = 36;
        weight_rom[1634] = 5;
        weight_rom[1635] = 41;
        weight_rom[1636] = 37;
        weight_rom[1637] = 34;
        weight_rom[1638] = 30;
        weight_rom[1639] = 32;
        weight_rom[1640] = 50;
        weight_rom[1641] = 46;
        weight_rom[1642] = 36;
        weight_rom[1643] = 19;
        weight_rom[1644] = 16;
        weight_rom[1645] = 8;
        weight_rom[1646] = -3;
        weight_rom[1647] = 17;
        weight_rom[1648] = 24;
        weight_rom[1649] = 25;
        weight_rom[1650] = 1;
        weight_rom[1651] = 1;
        weight_rom[1652] = 1;
        weight_rom[1653] = 0;
        weight_rom[1654] = -13;
        weight_rom[1655] = 0;
        weight_rom[1656] = 0;
        weight_rom[1657] = 38;
        weight_rom[1658] = 32;
        weight_rom[1659] = 23;
        weight_rom[1660] = 31;
        weight_rom[1661] = 29;
        weight_rom[1662] = 45;
        weight_rom[1663] = 19;
        weight_rom[1664] = 32;
        weight_rom[1665] = 33;
        weight_rom[1666] = 21;
        weight_rom[1667] = 21;
        weight_rom[1668] = 18;
        weight_rom[1669] = 21;
        weight_rom[1670] = 16;
        weight_rom[1671] = 9;
        weight_rom[1672] = 16;
        weight_rom[1673] = 4;
        weight_rom[1674] = -5;
        weight_rom[1675] = -1;
        weight_rom[1676] = -30;
        weight_rom[1677] = 15;
        weight_rom[1678] = -1;
        weight_rom[1679] = 0;
        weight_rom[1680] = 1;
        weight_rom[1681] = 2;
        weight_rom[1682] = 22;
        weight_rom[1683] = 1;
        weight_rom[1684] = -13;
        weight_rom[1685] = -2;
        weight_rom[1686] = 39;
        weight_rom[1687] = 19;
        weight_rom[1688] = 1;
        weight_rom[1689] = 18;
        weight_rom[1690] = 25;
        weight_rom[1691] = 9;
        weight_rom[1692] = 16;
        weight_rom[1693] = 16;
        weight_rom[1694] = 17;
        weight_rom[1695] = 13;
        weight_rom[1696] = 4;
        weight_rom[1697] = 4;
        weight_rom[1698] = 13;
        weight_rom[1699] = -2;
        weight_rom[1700] = -3;
        weight_rom[1701] = -8;
        weight_rom[1702] = -7;
        weight_rom[1703] = -9;
        weight_rom[1704] = -6;
        weight_rom[1705] = -2;
        weight_rom[1706] = 39;
        weight_rom[1707] = -1;
        weight_rom[1708] = 1;
        weight_rom[1709] = -1;
        weight_rom[1710] = 0;
        weight_rom[1711] = 22;
        weight_rom[1712] = 17;
        weight_rom[1713] = 12;
        weight_rom[1714] = 0;
        weight_rom[1715] = 13;
        weight_rom[1716] = 0;
        weight_rom[1717] = 6;
        weight_rom[1718] = 7;
        weight_rom[1719] = 7;
        weight_rom[1720] = 12;
        weight_rom[1721] = 11;
        weight_rom[1722] = 11;
        weight_rom[1723] = 10;
        weight_rom[1724] = 11;
        weight_rom[1725] = 6;
        weight_rom[1726] = 6;
        weight_rom[1727] = 2;
        weight_rom[1728] = 7;
        weight_rom[1729] = 0;
        weight_rom[1730] = 2;
        weight_rom[1731] = 1;
        weight_rom[1732] = 3;
        weight_rom[1733] = 12;
        weight_rom[1734] = 36;
        weight_rom[1735] = 0;
        weight_rom[1736] = 1;
        weight_rom[1737] = -2;
        weight_rom[1738] = 15;
        weight_rom[1739] = 40;
        weight_rom[1740] = 4;
        weight_rom[1741] = -1;
        weight_rom[1742] = 5;
        weight_rom[1743] = 3;
        weight_rom[1744] = 1;
        weight_rom[1745] = 9;
        weight_rom[1746] = 0;
        weight_rom[1747] = 1;
        weight_rom[1748] = 3;
        weight_rom[1749] = 7;
        weight_rom[1750] = 4;
        weight_rom[1751] = 6;
        weight_rom[1752] = 2;
        weight_rom[1753] = -1;
        weight_rom[1754] = 2;
        weight_rom[1755] = 0;
        weight_rom[1756] = -1;
        weight_rom[1757] = 0;
        weight_rom[1758] = -7;
        weight_rom[1759] = 0;
        weight_rom[1760] = 20;
        weight_rom[1761] = 13;
        weight_rom[1762] = 3;
        weight_rom[1763] = -4;
        weight_rom[1764] = 0;
        weight_rom[1765] = 30;
        weight_rom[1766] = 3;
        weight_rom[1767] = 4;
        weight_rom[1768] = 16;
        weight_rom[1769] = 5;
        weight_rom[1770] = 1;
        weight_rom[1771] = -10;
        weight_rom[1772] = 9;
        weight_rom[1773] = -9;
        weight_rom[1774] = 1;
        weight_rom[1775] = -4;
        weight_rom[1776] = -1;
        weight_rom[1777] = 1;
        weight_rom[1778] = 4;
        weight_rom[1779] = 3;
        weight_rom[1780] = -2;
        weight_rom[1781] = -3;
        weight_rom[1782] = -2;
        weight_rom[1783] = -4;
        weight_rom[1784] = -2;
        weight_rom[1785] = 0;
        weight_rom[1786] = 2;
        weight_rom[1787] = -5;
        weight_rom[1788] = 23;
        weight_rom[1789] = 28;
        weight_rom[1790] = 14;
        weight_rom[1791] = -32;
        weight_rom[1792] = 12;
        weight_rom[1793] = 14;
        weight_rom[1794] = 19;
        weight_rom[1795] = 11;
        weight_rom[1796] = 23;
        weight_rom[1797] = -3;
        weight_rom[1798] = 7;
        weight_rom[1799] = 2;
        weight_rom[1800] = -7;
        weight_rom[1801] = -4;
        weight_rom[1802] = 1;
        weight_rom[1803] = -3;
        weight_rom[1804] = 1;
        weight_rom[1805] = 6;
        weight_rom[1806] = 9;
        weight_rom[1807] = 1;
        weight_rom[1808] = -3;
        weight_rom[1809] = -1;
        weight_rom[1810] = -1;
        weight_rom[1811] = 2;
        weight_rom[1812] = 5;
        weight_rom[1813] = 0;
        weight_rom[1814] = 2;
        weight_rom[1815] = -1;
        weight_rom[1816] = 12;
        weight_rom[1817] = 23;
        weight_rom[1818] = 34;
        weight_rom[1819] = 29;
        weight_rom[1820] = 0;
        weight_rom[1821] = 25;
        weight_rom[1822] = -9;
        weight_rom[1823] = 21;
        weight_rom[1824] = 27;
        weight_rom[1825] = 0;
        weight_rom[1826] = 1;
        weight_rom[1827] = 3;
        weight_rom[1828] = -3;
        weight_rom[1829] = 3;
        weight_rom[1830] = -6;
        weight_rom[1831] = -4;
        weight_rom[1832] = -10;
        weight_rom[1833] = -2;
        weight_rom[1834] = 8;
        weight_rom[1835] = 1;
        weight_rom[1836] = -7;
        weight_rom[1837] = -4;
        weight_rom[1838] = -2;
        weight_rom[1839] = -3;
        weight_rom[1840] = -3;
        weight_rom[1841] = -8;
        weight_rom[1842] = 8;
        weight_rom[1843] = 2;
        weight_rom[1844] = 14;
        weight_rom[1845] = 34;
        weight_rom[1846] = 16;
        weight_rom[1847] = -9;
        weight_rom[1848] = 10;
        weight_rom[1849] = 7;
        weight_rom[1850] = -28;
        weight_rom[1851] = 14;
        weight_rom[1852] = 3;
        weight_rom[1853] = 15;
        weight_rom[1854] = 11;
        weight_rom[1855] = 5;
        weight_rom[1856] = -7;
        weight_rom[1857] = -10;
        weight_rom[1858] = -14;
        weight_rom[1859] = -14;
        weight_rom[1860] = -18;
        weight_rom[1861] = -19;
        weight_rom[1862] = 5;
        weight_rom[1863] = 3;
        weight_rom[1864] = -2;
        weight_rom[1865] = -10;
        weight_rom[1866] = -7;
        weight_rom[1867] = -12;
        weight_rom[1868] = -11;
        weight_rom[1869] = 2;
        weight_rom[1870] = -11;
        weight_rom[1871] = 1;
        weight_rom[1872] = 31;
        weight_rom[1873] = 48;
        weight_rom[1874] = 41;
        weight_rom[1875] = 17;
        weight_rom[1876] = 15;
        weight_rom[1877] = -12;
        weight_rom[1878] = 4;
        weight_rom[1879] = 5;
        weight_rom[1880] = 5;
        weight_rom[1881] = -3;
        weight_rom[1882] = -7;
        weight_rom[1883] = -15;
        weight_rom[1884] = -16;
        weight_rom[1885] = -18;
        weight_rom[1886] = -18;
        weight_rom[1887] = -16;
        weight_rom[1888] = -21;
        weight_rom[1889] = -13;
        weight_rom[1890] = 16;
        weight_rom[1891] = 7;
        weight_rom[1892] = -7;
        weight_rom[1893] = -7;
        weight_rom[1894] = -5;
        weight_rom[1895] = -3;
        weight_rom[1896] = -6;
        weight_rom[1897] = -13;
        weight_rom[1898] = -7;
        weight_rom[1899] = 1;
        weight_rom[1900] = 25;
        weight_rom[1901] = 50;
        weight_rom[1902] = 50;
        weight_rom[1903] = -25;
        weight_rom[1904] = 12;
        weight_rom[1905] = -11;
        weight_rom[1906] = -37;
        weight_rom[1907] = 1;
        weight_rom[1908] = -3;
        weight_rom[1909] = -8;
        weight_rom[1910] = -31;
        weight_rom[1911] = -21;
        weight_rom[1912] = -17;
        weight_rom[1913] = -12;
        weight_rom[1914] = -6;
        weight_rom[1915] = -10;
        weight_rom[1916] = -14;
        weight_rom[1917] = -5;
        weight_rom[1918] = 33;
        weight_rom[1919] = 14;
        weight_rom[1920] = -2;
        weight_rom[1921] = -3;
        weight_rom[1922] = 6;
        weight_rom[1923] = 6;
        weight_rom[1924] = 5;
        weight_rom[1925] = -2;
        weight_rom[1926] = -23;
        weight_rom[1927] = -21;
        weight_rom[1928] = -29;
        weight_rom[1929] = 29;
        weight_rom[1930] = 73;
        weight_rom[1931] = -22;
        weight_rom[1932] = 1;
        weight_rom[1933] = -11;
        weight_rom[1934] = -13;
        weight_rom[1935] = -17;
        weight_rom[1936] = -14;
        weight_rom[1937] = -37;
        weight_rom[1938] = -24;
        weight_rom[1939] = -20;
        weight_rom[1940] = -4;
        weight_rom[1941] = -4;
        weight_rom[1942] = -16;
        weight_rom[1943] = -9;
        weight_rom[1944] = -5;
        weight_rom[1945] = 10;
        weight_rom[1946] = 40;
        weight_rom[1947] = 10;
        weight_rom[1948] = -3;
        weight_rom[1949] = 1;
        weight_rom[1950] = 11;
        weight_rom[1951] = 4;
        weight_rom[1952] = -6;
        weight_rom[1953] = -15;
        weight_rom[1954] = -24;
        weight_rom[1955] = -23;
        weight_rom[1956] = -26;
        weight_rom[1957] = 27;
        weight_rom[1958] = 59;
        weight_rom[1959] = 0;
        weight_rom[1960] = -2;
        weight_rom[1961] = 1;
        weight_rom[1962] = -3;
        weight_rom[1963] = -9;
        weight_rom[1964] = -52;
        weight_rom[1965] = -39;
        weight_rom[1966] = -20;
        weight_rom[1967] = -6;
        weight_rom[1968] = -4;
        weight_rom[1969] = -8;
        weight_rom[1970] = -9;
        weight_rom[1971] = -4;
        weight_rom[1972] = -1;
        weight_rom[1973] = 19;
        weight_rom[1974] = 38;
        weight_rom[1975] = 14;
        weight_rom[1976] = -6;
        weight_rom[1977] = 4;
        weight_rom[1978] = 6;
        weight_rom[1979] = -6;
        weight_rom[1980] = -12;
        weight_rom[1981] = -10;
        weight_rom[1982] = -24;
        weight_rom[1983] = -26;
        weight_rom[1984] = -37;
        weight_rom[1985] = 1;
        weight_rom[1986] = 59;
        weight_rom[1987] = 1;
        weight_rom[1988] = -1;
        weight_rom[1989] = 22;
        weight_rom[1990] = 15;
        weight_rom[1991] = 12;
        weight_rom[1992] = -5;
        weight_rom[1993] = -18;
        weight_rom[1994] = -18;
        weight_rom[1995] = -11;
        weight_rom[1996] = -6;
        weight_rom[1997] = -8;
        weight_rom[1998] = -5;
        weight_rom[1999] = -7;
        weight_rom[2000] = 2;
        weight_rom[2001] = 33;
        weight_rom[2002] = 30;
        weight_rom[2003] = 9;
        weight_rom[2004] = -6;
        weight_rom[2005] = -5;
        weight_rom[2006] = -5;
        weight_rom[2007] = -5;
        weight_rom[2008] = -17;
        weight_rom[2009] = -16;
        weight_rom[2010] = -14;
        weight_rom[2011] = -21;
        weight_rom[2012] = 3;
        weight_rom[2013] = 33;
        weight_rom[2014] = 48;
        weight_rom[2015] = 25;
        weight_rom[2016] = 1;
        weight_rom[2017] = 0;
        weight_rom[2018] = 64;
        weight_rom[2019] = 51;
        weight_rom[2020] = 22;
        weight_rom[2021] = 6;
        weight_rom[2022] = 1;
        weight_rom[2023] = -3;
        weight_rom[2024] = -16;
        weight_rom[2025] = -3;
        weight_rom[2026] = -4;
        weight_rom[2027] = -1;
        weight_rom[2028] = 15;
        weight_rom[2029] = 32;
        weight_rom[2030] = 30;
        weight_rom[2031] = -2;
        weight_rom[2032] = -7;
        weight_rom[2033] = -2;
        weight_rom[2034] = -10;
        weight_rom[2035] = -10;
        weight_rom[2036] = -10;
        weight_rom[2037] = 1;
        weight_rom[2038] = 1;
        weight_rom[2039] = 6;
        weight_rom[2040] = 18;
        weight_rom[2041] = 77;
        weight_rom[2042] = 69;
        weight_rom[2043] = 46;
        weight_rom[2044] = -2;
        weight_rom[2045] = 18;
        weight_rom[2046] = 12;
        weight_rom[2047] = 39;
        weight_rom[2048] = 31;
        weight_rom[2049] = 5;
        weight_rom[2050] = 7;
        weight_rom[2051] = -2;
        weight_rom[2052] = -6;
        weight_rom[2053] = -4;
        weight_rom[2054] = 1;
        weight_rom[2055] = 2;
        weight_rom[2056] = 21;
        weight_rom[2057] = 23;
        weight_rom[2058] = 17;
        weight_rom[2059] = -5;
        weight_rom[2060] = -3;
        weight_rom[2061] = -3;
        weight_rom[2062] = -6;
        weight_rom[2063] = 0;
        weight_rom[2064] = -2;
        weight_rom[2065] = 2;
        weight_rom[2066] = -5;
        weight_rom[2067] = 6;
        weight_rom[2068] = 0;
        weight_rom[2069] = 69;
        weight_rom[2070] = 80;
        weight_rom[2071] = 1;
        weight_rom[2072] = 1;
        weight_rom[2073] = 17;
        weight_rom[2074] = 100;
        weight_rom[2075] = 35;
        weight_rom[2076] = 9;
        weight_rom[2077] = 13;
        weight_rom[2078] = 9;
        weight_rom[2079] = -5;
        weight_rom[2080] = 2;
        weight_rom[2081] = -3;
        weight_rom[2082] = 4;
        weight_rom[2083] = 5;
        weight_rom[2084] = 17;
        weight_rom[2085] = 21;
        weight_rom[2086] = 12;
        weight_rom[2087] = 1;
        weight_rom[2088] = 7;
        weight_rom[2089] = 5;
        weight_rom[2090] = 8;
        weight_rom[2091] = 10;
        weight_rom[2092] = 10;
        weight_rom[2093] = 8;
        weight_rom[2094] = 22;
        weight_rom[2095] = 19;
        weight_rom[2096] = 45;
        weight_rom[2097] = 81;
        weight_rom[2098] = 35;
        weight_rom[2099] = 30;
        weight_rom[2100] = 1;
        weight_rom[2101] = 20;
        weight_rom[2102] = -5;
        weight_rom[2103] = 37;
        weight_rom[2104] = 9;
        weight_rom[2105] = 10;
        weight_rom[2106] = 3;
        weight_rom[2107] = 11;
        weight_rom[2108] = 2;
        weight_rom[2109] = 11;
        weight_rom[2110] = 11;
        weight_rom[2111] = -1;
        weight_rom[2112] = 1;
        weight_rom[2113] = 10;
        weight_rom[2114] = 11;
        weight_rom[2115] = 12;
        weight_rom[2116] = 11;
        weight_rom[2117] = 13;
        weight_rom[2118] = 11;
        weight_rom[2119] = 6;
        weight_rom[2120] = 9;
        weight_rom[2121] = 10;
        weight_rom[2122] = 15;
        weight_rom[2123] = 18;
        weight_rom[2124] = 24;
        weight_rom[2125] = 68;
        weight_rom[2126] = 48;
        weight_rom[2127] = 20;
        weight_rom[2128] = 0;
        weight_rom[2129] = -11;
        weight_rom[2130] = -1;
        weight_rom[2131] = 40;
        weight_rom[2132] = 27;
        weight_rom[2133] = 12;
        weight_rom[2134] = 16;
        weight_rom[2135] = 12;
        weight_rom[2136] = 14;
        weight_rom[2137] = 14;
        weight_rom[2138] = 11;
        weight_rom[2139] = 7;
        weight_rom[2140] = -5;
        weight_rom[2141] = -7;
        weight_rom[2142] = 4;
        weight_rom[2143] = 5;
        weight_rom[2144] = 5;
        weight_rom[2145] = 9;
        weight_rom[2146] = 12;
        weight_rom[2147] = 5;
        weight_rom[2148] = 14;
        weight_rom[2149] = 11;
        weight_rom[2150] = 5;
        weight_rom[2151] = 28;
        weight_rom[2152] = 55;
        weight_rom[2153] = 25;
        weight_rom[2154] = 13;
        weight_rom[2155] = -1;
        weight_rom[2156] = -2;
        weight_rom[2157] = -1;
        weight_rom[2158] = 46;
        weight_rom[2159] = 63;
        weight_rom[2160] = 5;
        weight_rom[2161] = 7;
        weight_rom[2162] = 10;
        weight_rom[2163] = 10;
        weight_rom[2164] = 11;
        weight_rom[2165] = 7;
        weight_rom[2166] = 3;
        weight_rom[2167] = -3;
        weight_rom[2168] = -7;
        weight_rom[2169] = -1;
        weight_rom[2170] = -1;
        weight_rom[2171] = -2;
        weight_rom[2172] = 0;
        weight_rom[2173] = 6;
        weight_rom[2174] = 6;
        weight_rom[2175] = 14;
        weight_rom[2176] = 5;
        weight_rom[2177] = 6;
        weight_rom[2178] = 12;
        weight_rom[2179] = 30;
        weight_rom[2180] = 31;
        weight_rom[2181] = 22;
        weight_rom[2182] = 4;
        weight_rom[2183] = -2;
        weight_rom[2184] = 2;
        weight_rom[2185] = -1;
        weight_rom[2186] = 69;
        weight_rom[2187] = 38;
        weight_rom[2188] = 27;
        weight_rom[2189] = 11;
        weight_rom[2190] = 13;
        weight_rom[2191] = 10;
        weight_rom[2192] = 2;
        weight_rom[2193] = 3;
        weight_rom[2194] = -1;
        weight_rom[2195] = 5;
        weight_rom[2196] = -2;
        weight_rom[2197] = -5;
        weight_rom[2198] = 0;
        weight_rom[2199] = 2;
        weight_rom[2200] = -4;
        weight_rom[2201] = 2;
        weight_rom[2202] = 4;
        weight_rom[2203] = 6;
        weight_rom[2204] = 13;
        weight_rom[2205] = 6;
        weight_rom[2206] = 13;
        weight_rom[2207] = 13;
        weight_rom[2208] = 25;
        weight_rom[2209] = -2;
        weight_rom[2210] = 19;
        weight_rom[2211] = -1;
        weight_rom[2212] = -1;
        weight_rom[2213] = 1;
        weight_rom[2214] = 49;
        weight_rom[2215] = 45;
        weight_rom[2216] = 38;
        weight_rom[2217] = 7;
        weight_rom[2218] = 13;
        weight_rom[2219] = 0;
        weight_rom[2220] = 8;
        weight_rom[2221] = 10;
        weight_rom[2222] = 1;
        weight_rom[2223] = 2;
        weight_rom[2224] = 7;
        weight_rom[2225] = 6;
        weight_rom[2226] = 4;
        weight_rom[2227] = 4;
        weight_rom[2228] = 7;
        weight_rom[2229] = -5;
        weight_rom[2230] = 3;
        weight_rom[2231] = 11;
        weight_rom[2232] = 19;
        weight_rom[2233] = 7;
        weight_rom[2234] = 20;
        weight_rom[2235] = 11;
        weight_rom[2236] = 0;
        weight_rom[2237] = 3;
        weight_rom[2238] = 13;
        weight_rom[2239] = -1;
        weight_rom[2240] = 1;
        weight_rom[2241] = 1;
        weight_rom[2242] = 25;
        weight_rom[2243] = 21;
        weight_rom[2244] = 9;
        weight_rom[2245] = 0;
        weight_rom[2246] = 5;
        weight_rom[2247] = 4;
        weight_rom[2248] = 1;
        weight_rom[2249] = 6;
        weight_rom[2250] = -2;
        weight_rom[2251] = 13;
        weight_rom[2252] = 12;
        weight_rom[2253] = 7;
        weight_rom[2254] = 14;
        weight_rom[2255] = 10;
        weight_rom[2256] = 12;
        weight_rom[2257] = 5;
        weight_rom[2258] = 3;
        weight_rom[2259] = -6;
        weight_rom[2260] = -18;
        weight_rom[2261] = 0;
        weight_rom[2262] = 1;
        weight_rom[2263] = -18;
        weight_rom[2264] = 24;
        weight_rom[2265] = 13;
        weight_rom[2266] = 0;
        weight_rom[2267] = 0;
        weight_rom[2268] = 0;
        weight_rom[2269] = 2;
        weight_rom[2270] = -1;
        weight_rom[2271] = -1;
        weight_rom[2272] = -14;
        weight_rom[2273] = -34;
        weight_rom[2274] = 6;
        weight_rom[2275] = -23;
        weight_rom[2276] = 8;
        weight_rom[2277] = -2;
        weight_rom[2278] = 3;
        weight_rom[2279] = -4;
        weight_rom[2280] = 7;
        weight_rom[2281] = -7;
        weight_rom[2282] = 9;
        weight_rom[2283] = -6;
        weight_rom[2284] = -1;
        weight_rom[2285] = 11;
        weight_rom[2286] = 2;
        weight_rom[2287] = 0;
        weight_rom[2288] = -12;
        weight_rom[2289] = -36;
        weight_rom[2290] = 2;
        weight_rom[2291] = -10;
        weight_rom[2292] = 20;
        weight_rom[2293] = -1;
        weight_rom[2294] = 1;
        weight_rom[2295] = -1;
        weight_rom[2296] = 0;
        weight_rom[2297] = -1;
        weight_rom[2298] = -1;
        weight_rom[2299] = 1;
        weight_rom[2300] = -37;
        weight_rom[2301] = -47;
        weight_rom[2302] = -13;
        weight_rom[2303] = -17;
        weight_rom[2304] = -15;
        weight_rom[2305] = 6;
        weight_rom[2306] = -4;
        weight_rom[2307] = 2;
        weight_rom[2308] = 13;
        weight_rom[2309] = 7;
        weight_rom[2310] = -1;
        weight_rom[2311] = 2;
        weight_rom[2312] = -1;
        weight_rom[2313] = 12;
        weight_rom[2314] = 11;
        weight_rom[2315] = 6;
        weight_rom[2316] = 13;
        weight_rom[2317] = -23;
        weight_rom[2318] = -14;
        weight_rom[2319] = -3;
        weight_rom[2320] = -2;
        weight_rom[2321] = -1;
        weight_rom[2322] = -1;
        weight_rom[2323] = -1;
        weight_rom[2324] = 0;
        weight_rom[2325] = 1;
        weight_rom[2326] = 0;
        weight_rom[2327] = 1;
        weight_rom[2328] = 1;
        weight_rom[2329] = 3;
        weight_rom[2330] = 3;
        weight_rom[2331] = 10;
        weight_rom[2332] = 1;
        weight_rom[2333] = -7;
        weight_rom[2334] = 3;
        weight_rom[2335] = 13;
        weight_rom[2336] = 30;
        weight_rom[2337] = 29;
        weight_rom[2338] = 17;
        weight_rom[2339] = 31;
        weight_rom[2340] = 19;
        weight_rom[2341] = 67;
        weight_rom[2342] = -24;
        weight_rom[2343] = 29;
        weight_rom[2344] = -11;
        weight_rom[2345] = -9;
        weight_rom[2346] = -26;
        weight_rom[2347] = -2;
        weight_rom[2348] = 0;
        weight_rom[2349] = -1;
        weight_rom[2350] = 0;
        weight_rom[2351] = -1;
        weight_rom[2352] = 127;
        weight_rom[2353] = 63;
        weight_rom[2354] = 20;
        weight_rom[2355] = -127;
        weight_rom[2356] = -29;
        weight_rom[2357] = -67;
        weight_rom[2358] = 29;
        weight_rom[2359] = -34;
        weight_rom[2360] = 36;
        weight_rom[2361] = -51;
        weight_rom[2362] = -10;
        weight_rom[2363] = 51;
        weight_rom[2364] = -19;
        weight_rom[2365] = -66;
        weight_rom[2366] = 54;
        weight_rom[2367] = 0;
        weight_rom[2368] = 43;
        weight_rom[2369] = -86;
        weight_rom[2370] = -59;
        weight_rom[2371] = -3;
        weight_rom[2372] = 0;
        weight_rom[2373] = -96;
        weight_rom[2374] = 57;
        weight_rom[2375] = -34;
        weight_rom[2376] = 75;
        weight_rom[2377] = -95;
        weight_rom[2378] = -23;
        weight_rom[2379] = -16;
        weight_rom[2380] = 18;
        weight_rom[2381] = 11;
        weight_rom[2382] = 59;
        weight_rom[2383] = -16;
        weight_rom[2384] = -61;
        weight_rom[2385] = 127;
        weight_rom[2386] = -94;
        weight_rom[2387] = -42;
        weight_rom[2388] = 8;
        weight_rom[2389] = -32;
        weight_rom[2390] = 65;
        weight_rom[2391] = -40;
        weight_rom[2392] = -11;
        weight_rom[2393] = -46;
        weight_rom[2394] = -35;
    end

    // 主状态机和MAC单元
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            valid <= 0;
            digit_out <= 0;
            neuron_idx <= 0;
            input_idx <= 0;
            accumulator <= 0;
            layer1_done <= 0;
        end else begin
            case (state)
                IDLE: begin
                    valid <= 0;
                    if (start) begin
                        state <= LAYER1;
                        neuron_idx <= 0;
                        input_idx <= 0;
                        layer1_done <= 0;
                        accumulator <= $signed({{16{weight_rom[2352][7]}}, weight_rom[2352]});
                    end
                end

                LAYER1: begin
                    // Layer1 MAC: acc += weight * input
                    if (input_idx < 784) begin
                        accumulator <= accumulator + ($signed({{16{weight_rom[neuron_idx * 784 + input_idx][7]}}, weight_rom[neuron_idx * 784 + input_idx]}) * $signed({23'b0, image_in[input_idx]}));
                        input_idx <= input_idx + 1;
                    end else begin
                        // ReLU并存储
                        layer1_out[neuron_idx] <= (accumulator[23] == 1'b1) ? 24'b0 : accumulator;

                        if (neuron_idx == 2) begin
                            // Layer1完成
                            state <= LAYER2;
                            neuron_idx <= 0;
                            input_idx <= 0;
                            accumulator <= $signed({{16{weight_rom[2385][7]}}, weight_rom[2385]});
                        end else begin
                            // 下一个神经元
                            neuron_idx <= neuron_idx + 1;
                            input_idx <= 0;
                            accumulator <= $signed({{16{weight_rom[2352 + neuron_idx + 1][7]}}, weight_rom[2352 + neuron_idx + 1]});
                        end
                    end
                end

                LAYER2: begin
                    // Layer2 MAC: acc += (weight * layer1_out) >> 7
                    if (input_idx < 3) begin
                        accumulator <= accumulator + (($signed({{16{weight_rom[2355 + neuron_idx * 3 + input_idx][7]}}, weight_rom[2355 + neuron_idx * 3 + input_idx]}) * layer1_out[input_idx]) >>> 7);
                        input_idx <= input_idx + 1;
                    end else begin
                        // 存储输出
                        layer2_out[neuron_idx] <= accumulator;

                        if (neuron_idx == 9) begin
                            // Layer2完成，进入argmax
                            state <= ARGMAX;
                            neuron_idx <= 0;
                            input_idx <= 0;
                            max_idx <= 0;
                            max_val <= layer2_out[0];
                        end else begin
                            // 下一个神经元
                            neuron_idx <= neuron_idx + 1;
                            input_idx <= 0;
                            accumulator <= $signed({{16{weight_rom[2385 + neuron_idx + 1][7]}}, weight_rom[2385 + neuron_idx + 1]});
                        end
                    end
                end

                ARGMAX: begin
                    // 串行比较查找最大值
                    if (input_idx == 0) begin
                        // 初始化已在LAYER2完成
                        input_idx <= 1;
                    end else if (input_idx < 10) begin
                        if (layer2_out[input_idx] > max_val) begin
                            max_val <= layer2_out[input_idx];
                            max_idx <= input_idx[3:0];
                        end
                        input_idx <= input_idx + 1;
                    end else begin
                        // 完成
                        digit_out <= max_idx;
                        valid <= 1;
                        state <= IDLE;
                        input_idx <= 0;
                    end
                end

                default: state <= IDLE;
            endcase
        end
    end

endmodule
