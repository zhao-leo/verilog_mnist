// MNIST手写数字识别模型 - Int8量化版本（串行计算架构）
// 架构优化：使用单个MAC单元串行计算，大幅减少逻辑门数量
// 输入: 28x28二值图像 (784位)
// 输出: 预测数字 (0-9)
// 时钟周期: ~13000 (Layer1: 16×784=12544 + Layer2: 10×16=160 + 其他)
// ROM布局: Layer1权重[0:12543] + Layer1偏置[12544:12559] +
//          Layer2权重[12560:12719] + Layer2偏置[12720:12729]

module mnist_model(
    input wire clk,
    input wire rst,
    input wire [783:0] image_in,  // 28*28 = 784位输入
    input wire start,
    output reg [3:0] digit_out,   // 输出数字 0-9
    output reg valid
);

    // 状态机
    localparam IDLE = 3'd0;
    localparam LAYER1_COMPUTE = 3'd1;
    localparam LAYER1_ACTIVATE = 3'd2;
    localparam LAYER2_COMPUTE = 3'd3;
    localparam ARGMAX = 3'd4;
    localparam DONE = 3'd5;

    reg [2:0] state;
    reg [4:0] neuron_idx;       // 当前神经元索引 (0-15 for layer1, 0-9 for layer2)
    reg [9:0] input_idx;        // 当前输入索引 (0-783 for layer1, 0-15 for layer2)

    // MAC单元
    reg signed [31:0] accumulator; // 累加器

    // 层输出存储
    reg signed [31:0] layer1_out [0:15];
    reg signed [31:0] layer2_out [0:9];

    // ROM: 存储所有权重和偏置 (12730个Int8参数)
    reg signed [7:0] weight_rom [0:12729];

    // 初始化ROM
    initial begin
        weight_rom[0] = 2;
        weight_rom[1] = 1;
        weight_rom[2] = -4;
        weight_rom[3] = 4;
        weight_rom[4] = -1;
        weight_rom[5] = -1;
        weight_rom[6] = -3;
        weight_rom[7] = 0;
        weight_rom[8] = -1;
        weight_rom[9] = 0;
        weight_rom[10] = 2;
        weight_rom[11] = 3;
        weight_rom[12] = -3;
        weight_rom[13] = 3;
        weight_rom[14] = 1;
        weight_rom[15] = 3;
        weight_rom[16] = -1;
        weight_rom[17] = 3;
        weight_rom[18] = 4;
        weight_rom[19] = 0;
        weight_rom[20] = 3;
        weight_rom[21] = 3;
        weight_rom[22] = 1;
        weight_rom[23] = 0;
        weight_rom[24] = 4;
        weight_rom[25] = -4;
        weight_rom[26] = 2;
        weight_rom[27] = -2;
        weight_rom[28] = -2;
        weight_rom[29] = 0;
        weight_rom[30] = 4;
        weight_rom[31] = -1;
        weight_rom[32] = 0;
        weight_rom[33] = -1;
        weight_rom[34] = -2;
        weight_rom[35] = -4;
        weight_rom[36] = -6;
        weight_rom[37] = -3;
        weight_rom[38] = -11;
        weight_rom[39] = -15;
        weight_rom[40] = -25;
        weight_rom[41] = -25;
        weight_rom[42] = -9;
        weight_rom[43] = 4;
        weight_rom[44] = -14;
        weight_rom[45] = -11;
        weight_rom[46] = -22;
        weight_rom[47] = -20;
        weight_rom[48] = -20;
        weight_rom[49] = -11;
        weight_rom[50] = -8;
        weight_rom[51] = -16;
        weight_rom[52] = 4;
        weight_rom[53] = 3;
        weight_rom[54] = 0;
        weight_rom[55] = 0;
        weight_rom[56] = 2;
        weight_rom[57] = 1;
        weight_rom[58] = 1;
        weight_rom[59] = 2;
        weight_rom[60] = -10;
        weight_rom[61] = 4;
        weight_rom[62] = -14;
        weight_rom[63] = -12;
        weight_rom[64] = -22;
        weight_rom[65] = -38;
        weight_rom[66] = -30;
        weight_rom[67] = -38;
        weight_rom[68] = -29;
        weight_rom[69] = 6;
        weight_rom[70] = -24;
        weight_rom[71] = 5;
        weight_rom[72] = 4;
        weight_rom[73] = 16;
        weight_rom[74] = 10;
        weight_rom[75] = 5;
        weight_rom[76] = -17;
        weight_rom[77] = -9;
        weight_rom[78] = -19;
        weight_rom[79] = -25;
        weight_rom[80] = -26;
        weight_rom[81] = -21;
        weight_rom[82] = -4;
        weight_rom[83] = 4;
        weight_rom[84] = -4;
        weight_rom[85] = -2;
        weight_rom[86] = -8;
        weight_rom[87] = -3;
        weight_rom[88] = 4;
        weight_rom[89] = -4;
        weight_rom[90] = -6;
        weight_rom[91] = -25;
        weight_rom[92] = -10;
        weight_rom[93] = 5;
        weight_rom[94] = -1;
        weight_rom[95] = -21;
        weight_rom[96] = -7;
        weight_rom[97] = -4;
        weight_rom[98] = -7;
        weight_rom[99] = 13;
        weight_rom[100] = 15;
        weight_rom[101] = 5;
        weight_rom[102] = 12;
        weight_rom[103] = 7;
        weight_rom[104] = 19;
        weight_rom[105] = 12;
        weight_rom[106] = 1;
        weight_rom[107] = -1;
        weight_rom[108] = -10;
        weight_rom[109] = 20;
        weight_rom[110] = 0;
        weight_rom[111] = 0;
        weight_rom[112] = 4;
        weight_rom[113] = 0;
        weight_rom[114] = 14;
        weight_rom[115] = 4;
        weight_rom[116] = -1;
        weight_rom[117] = -14;
        weight_rom[118] = -28;
        weight_rom[119] = -12;
        weight_rom[120] = -8;
        weight_rom[121] = -9;
        weight_rom[122] = 2;
        weight_rom[123] = 6;
        weight_rom[124] = 1;
        weight_rom[125] = 16;
        weight_rom[126] = 20;
        weight_rom[127] = 18;
        weight_rom[128] = 19;
        weight_rom[129] = 4;
        weight_rom[130] = 21;
        weight_rom[131] = 7;
        weight_rom[132] = 10;
        weight_rom[133] = 15;
        weight_rom[134] = -13;
        weight_rom[135] = 7;
        weight_rom[136] = 13;
        weight_rom[137] = 17;
        weight_rom[138] = 10;
        weight_rom[139] = 4;
        weight_rom[140] = 4;
        weight_rom[141] = 2;
        weight_rom[142] = -3;
        weight_rom[143] = 12;
        weight_rom[144] = -25;
        weight_rom[145] = 16;
        weight_rom[146] = -5;
        weight_rom[147] = -6;
        weight_rom[148] = -5;
        weight_rom[149] = -1;
        weight_rom[150] = -7;
        weight_rom[151] = 2;
        weight_rom[152] = -8;
        weight_rom[153] = -9;
        weight_rom[154] = -1;
        weight_rom[155] = -7;
        weight_rom[156] = -4;
        weight_rom[157] = -14;
        weight_rom[158] = -12;
        weight_rom[159] = -4;
        weight_rom[160] = -3;
        weight_rom[161] = -4;
        weight_rom[162] = -2;
        weight_rom[163] = 6;
        weight_rom[164] = 1;
        weight_rom[165] = 14;
        weight_rom[166] = 6;
        weight_rom[167] = -3;
        weight_rom[168] = -1;
        weight_rom[169] = 4;
        weight_rom[170] = 14;
        weight_rom[171] = 1;
        weight_rom[172] = 2;
        weight_rom[173] = -4;
        weight_rom[174] = 0;
        weight_rom[175] = -12;
        weight_rom[176] = -11;
        weight_rom[177] = 1;
        weight_rom[178] = 11;
        weight_rom[179] = 12;
        weight_rom[180] = 1;
        weight_rom[181] = -5;
        weight_rom[182] = -3;
        weight_rom[183] = -3;
        weight_rom[184] = -3;
        weight_rom[185] = -7;
        weight_rom[186] = 1;
        weight_rom[187] = 4;
        weight_rom[188] = 7;
        weight_rom[189] = 5;
        weight_rom[190] = -8;
        weight_rom[191] = -2;
        weight_rom[192] = 33;
        weight_rom[193] = 28;
        weight_rom[194] = 11;
        weight_rom[195] = -2;
        weight_rom[196] = 1;
        weight_rom[197] = 3;
        weight_rom[198] = 9;
        weight_rom[199] = 9;
        weight_rom[200] = -17;
        weight_rom[201] = -10;
        weight_rom[202] = -6;
        weight_rom[203] = 9;
        weight_rom[204] = 3;
        weight_rom[205] = 6;
        weight_rom[206] = 15;
        weight_rom[207] = 12;
        weight_rom[208] = 9;
        weight_rom[209] = 1;
        weight_rom[210] = 10;
        weight_rom[211] = -1;
        weight_rom[212] = 2;
        weight_rom[213] = 9;
        weight_rom[214] = 12;
        weight_rom[215] = 15;
        weight_rom[216] = 15;
        weight_rom[217] = 14;
        weight_rom[218] = 8;
        weight_rom[219] = 14;
        weight_rom[220] = 6;
        weight_rom[221] = 16;
        weight_rom[222] = 2;
        weight_rom[223] = 0;
        weight_rom[224] = 10;
        weight_rom[225] = 11;
        weight_rom[226] = -2;
        weight_rom[227] = 10;
        weight_rom[228] = -9;
        weight_rom[229] = -3;
        weight_rom[230] = 4;
        weight_rom[231] = 12;
        weight_rom[232] = 6;
        weight_rom[233] = 5;
        weight_rom[234] = 13;
        weight_rom[235] = 22;
        weight_rom[236] = 24;
        weight_rom[237] = 22;
        weight_rom[238] = 21;
        weight_rom[239] = 12;
        weight_rom[240] = 7;
        weight_rom[241] = 14;
        weight_rom[242] = 14;
        weight_rom[243] = 15;
        weight_rom[244] = 16;
        weight_rom[245] = 20;
        weight_rom[246] = 22;
        weight_rom[247] = 23;
        weight_rom[248] = 27;
        weight_rom[249] = 41;
        weight_rom[250] = 40;
        weight_rom[251] = 1;
        weight_rom[252] = 13;
        weight_rom[253] = 15;
        weight_rom[254] = 7;
        weight_rom[255] = 12;
        weight_rom[256] = 4;
        weight_rom[257] = 3;
        weight_rom[258] = 3;
        weight_rom[259] = -3;
        weight_rom[260] = 11;
        weight_rom[261] = 9;
        weight_rom[262] = 4;
        weight_rom[263] = 28;
        weight_rom[264] = 33;
        weight_rom[265] = 19;
        weight_rom[266] = 22;
        weight_rom[267] = 19;
        weight_rom[268] = 10;
        weight_rom[269] = 5;
        weight_rom[270] = -1;
        weight_rom[271] = 3;
        weight_rom[272] = 10;
        weight_rom[273] = 27;
        weight_rom[274] = 21;
        weight_rom[275] = 11;
        weight_rom[276] = 49;
        weight_rom[277] = 70;
        weight_rom[278] = 28;
        weight_rom[279] = 14;
        weight_rom[280] = 16;
        weight_rom[281] = 19;
        weight_rom[282] = 2;
        weight_rom[283] = 10;
        weight_rom[284] = 5;
        weight_rom[285] = -3;
        weight_rom[286] = -7;
        weight_rom[287] = -3;
        weight_rom[288] = 0;
        weight_rom[289] = 5;
        weight_rom[290] = 17;
        weight_rom[291] = 19;
        weight_rom[292] = 30;
        weight_rom[293] = 34;
        weight_rom[294] = 45;
        weight_rom[295] = 26;
        weight_rom[296] = 22;
        weight_rom[297] = 2;
        weight_rom[298] = -2;
        weight_rom[299] = 0;
        weight_rom[300] = -6;
        weight_rom[301] = 7;
        weight_rom[302] = -3;
        weight_rom[303] = 14;
        weight_rom[304] = 34;
        weight_rom[305] = 81;
        weight_rom[306] = 48;
        weight_rom[307] = 17;
        weight_rom[308] = 18;
        weight_rom[309] = 15;
        weight_rom[310] = 30;
        weight_rom[311] = 6;
        weight_rom[312] = 22;
        weight_rom[313] = 0;
        weight_rom[314] = -2;
        weight_rom[315] = -4;
        weight_rom[316] = -18;
        weight_rom[317] = -11;
        weight_rom[318] = 2;
        weight_rom[319] = 6;
        weight_rom[320] = 10;
        weight_rom[321] = 24;
        weight_rom[322] = 30;
        weight_rom[323] = 30;
        weight_rom[324] = 15;
        weight_rom[325] = 3;
        weight_rom[326] = -1;
        weight_rom[327] = -25;
        weight_rom[328] = -32;
        weight_rom[329] = -37;
        weight_rom[330] = -30;
        weight_rom[331] = -24;
        weight_rom[332] = -19;
        weight_rom[333] = 44;
        weight_rom[334] = 31;
        weight_rom[335] = -2;
        weight_rom[336] = 9;
        weight_rom[337] = 13;
        weight_rom[338] = 19;
        weight_rom[339] = 17;
        weight_rom[340] = 19;
        weight_rom[341] = 4;
        weight_rom[342] = -12;
        weight_rom[343] = -14;
        weight_rom[344] = -15;
        weight_rom[345] = -20;
        weight_rom[346] = -21;
        weight_rom[347] = -19;
        weight_rom[348] = -32;
        weight_rom[349] = -17;
        weight_rom[350] = 26;
        weight_rom[351] = 26;
        weight_rom[352] = 7;
        weight_rom[353] = -6;
        weight_rom[354] = -3;
        weight_rom[355] = -30;
        weight_rom[356] = -34;
        weight_rom[357] = -53;
        weight_rom[358] = -65;
        weight_rom[359] = -63;
        weight_rom[360] = -71;
        weight_rom[361] = -16;
        weight_rom[362] = 14;
        weight_rom[363] = 2;
        weight_rom[364] = 4;
        weight_rom[365] = 3;
        weight_rom[366] = 27;
        weight_rom[367] = 5;
        weight_rom[368] = 11;
        weight_rom[369] = -17;
        weight_rom[370] = -16;
        weight_rom[371] = -16;
        weight_rom[372] = -24;
        weight_rom[373] = -24;
        weight_rom[374] = -45;
        weight_rom[375] = -50;
        weight_rom[376] = -34;
        weight_rom[377] = -6;
        weight_rom[378] = 21;
        weight_rom[379] = 15;
        weight_rom[380] = 3;
        weight_rom[381] = 3;
        weight_rom[382] = 0;
        weight_rom[383] = -10;
        weight_rom[384] = -22;
        weight_rom[385] = -49;
        weight_rom[386] = -54;
        weight_rom[387] = -66;
        weight_rom[388] = -44;
        weight_rom[389] = -24;
        weight_rom[390] = -26;
        weight_rom[391] = -10;
        weight_rom[392] = 0;
        weight_rom[393] = 3;
        weight_rom[394] = 21;
        weight_rom[395] = 8;
        weight_rom[396] = 1;
        weight_rom[397] = -12;
        weight_rom[398] = -19;
        weight_rom[399] = -28;
        weight_rom[400] = -37;
        weight_rom[401] = -38;
        weight_rom[402] = -28;
        weight_rom[403] = -51;
        weight_rom[404] = -37;
        weight_rom[405] = -2;
        weight_rom[406] = 34;
        weight_rom[407] = 9;
        weight_rom[408] = 6;
        weight_rom[409] = 2;
        weight_rom[410] = 6;
        weight_rom[411] = 7;
        weight_rom[412] = 3;
        weight_rom[413] = -17;
        weight_rom[414] = -24;
        weight_rom[415] = -29;
        weight_rom[416] = -44;
        weight_rom[417] = -23;
        weight_rom[418] = -6;
        weight_rom[419] = -3;
        weight_rom[420] = -1;
        weight_rom[421] = 12;
        weight_rom[422] = 28;
        weight_rom[423] = 1;
        weight_rom[424] = -15;
        weight_rom[425] = -25;
        weight_rom[426] = -3;
        weight_rom[427] = -27;
        weight_rom[428] = -29;
        weight_rom[429] = -30;
        weight_rom[430] = -25;
        weight_rom[431] = -32;
        weight_rom[432] = -20;
        weight_rom[433] = 0;
        weight_rom[434] = 13;
        weight_rom[435] = 10;
        weight_rom[436] = -9;
        weight_rom[437] = -6;
        weight_rom[438] = 18;
        weight_rom[439] = 2;
        weight_rom[440] = 12;
        weight_rom[441] = 1;
        weight_rom[442] = -8;
        weight_rom[443] = -15;
        weight_rom[444] = -13;
        weight_rom[445] = -30;
        weight_rom[446] = -7;
        weight_rom[447] = -3;
        weight_rom[448] = 1;
        weight_rom[449] = 1;
        weight_rom[450] = -2;
        weight_rom[451] = 4;
        weight_rom[452] = 5;
        weight_rom[453] = -9;
        weight_rom[454] = 3;
        weight_rom[455] = -15;
        weight_rom[456] = -23;
        weight_rom[457] = -20;
        weight_rom[458] = -25;
        weight_rom[459] = -28;
        weight_rom[460] = -12;
        weight_rom[461] = 8;
        weight_rom[462] = 1;
        weight_rom[463] = 4;
        weight_rom[464] = 3;
        weight_rom[465] = -2;
        weight_rom[466] = 5;
        weight_rom[467] = 16;
        weight_rom[468] = 5;
        weight_rom[469] = -3;
        weight_rom[470] = -4;
        weight_rom[471] = -31;
        weight_rom[472] = -25;
        weight_rom[473] = -16;
        weight_rom[474] = 5;
        weight_rom[475] = -11;
        weight_rom[476] = -4;
        weight_rom[477] = -5;
        weight_rom[478] = -23;
        weight_rom[479] = -1;
        weight_rom[480] = 18;
        weight_rom[481] = -2;
        weight_rom[482] = 9;
        weight_rom[483] = 4;
        weight_rom[484] = 2;
        weight_rom[485] = -6;
        weight_rom[486] = -16;
        weight_rom[487] = -24;
        weight_rom[488] = -17;
        weight_rom[489] = 3;
        weight_rom[490] = 13;
        weight_rom[491] = 12;
        weight_rom[492] = 6;
        weight_rom[493] = 9;
        weight_rom[494] = 5;
        weight_rom[495] = 3;
        weight_rom[496] = 11;
        weight_rom[497] = 1;
        weight_rom[498] = -15;
        weight_rom[499] = -16;
        weight_rom[500] = -13;
        weight_rom[501] = -22;
        weight_rom[502] = -2;
        weight_rom[503] = -1;
        weight_rom[504] = -3;
        weight_rom[505] = -5;
        weight_rom[506] = 1;
        weight_rom[507] = 10;
        weight_rom[508] = 23;
        weight_rom[509] = -1;
        weight_rom[510] = 4;
        weight_rom[511] = 10;
        weight_rom[512] = 14;
        weight_rom[513] = 6;
        weight_rom[514] = -18;
        weight_rom[515] = -10;
        weight_rom[516] = -17;
        weight_rom[517] = 15;
        weight_rom[518] = 25;
        weight_rom[519] = 13;
        weight_rom[520] = -5;
        weight_rom[521] = 6;
        weight_rom[522] = 11;
        weight_rom[523] = 11;
        weight_rom[524] = 6;
        weight_rom[525] = -4;
        weight_rom[526] = -9;
        weight_rom[527] = -22;
        weight_rom[528] = -38;
        weight_rom[529] = -32;
        weight_rom[530] = 3;
        weight_rom[531] = 14;
        weight_rom[532] = 0;
        weight_rom[533] = -5;
        weight_rom[534] = 14;
        weight_rom[535] = 3;
        weight_rom[536] = 11;
        weight_rom[537] = -9;
        weight_rom[538] = 1;
        weight_rom[539] = 13;
        weight_rom[540] = 20;
        weight_rom[541] = 18;
        weight_rom[542] = -7;
        weight_rom[543] = -8;
        weight_rom[544] = -3;
        weight_rom[545] = 13;
        weight_rom[546] = 21;
        weight_rom[547] = 15;
        weight_rom[548] = 9;
        weight_rom[549] = 6;
        weight_rom[550] = 5;
        weight_rom[551] = 11;
        weight_rom[552] = 1;
        weight_rom[553] = -13;
        weight_rom[554] = -20;
        weight_rom[555] = -20;
        weight_rom[556] = 1;
        weight_rom[557] = -7;
        weight_rom[558] = -11;
        weight_rom[559] = -2;
        weight_rom[560] = 3;
        weight_rom[561] = -18;
        weight_rom[562] = 5;
        weight_rom[563] = -3;
        weight_rom[564] = -25;
        weight_rom[565] = -13;
        weight_rom[566] = 3;
        weight_rom[567] = -6;
        weight_rom[568] = 10;
        weight_rom[569] = 5;
        weight_rom[570] = 1;
        weight_rom[571] = -1;
        weight_rom[572] = 1;
        weight_rom[573] = 4;
        weight_rom[574] = 15;
        weight_rom[575] = 6;
        weight_rom[576] = 7;
        weight_rom[577] = 11;
        weight_rom[578] = 3;
        weight_rom[579] = 5;
        weight_rom[580] = -11;
        weight_rom[581] = -20;
        weight_rom[582] = -17;
        weight_rom[583] = -16;
        weight_rom[584] = 5;
        weight_rom[585] = -6;
        weight_rom[586] = -6;
        weight_rom[587] = 3;
        weight_rom[588] = -4;
        weight_rom[589] = -14;
        weight_rom[590] = -17;
        weight_rom[591] = -12;
        weight_rom[592] = -3;
        weight_rom[593] = -1;
        weight_rom[594] = 2;
        weight_rom[595] = 3;
        weight_rom[596] = 2;
        weight_rom[597] = 5;
        weight_rom[598] = 3;
        weight_rom[599] = -2;
        weight_rom[600] = 3;
        weight_rom[601] = 4;
        weight_rom[602] = 1;
        weight_rom[603] = 3;
        weight_rom[604] = 1;
        weight_rom[605] = 1;
        weight_rom[606] = -3;
        weight_rom[607] = 1;
        weight_rom[608] = -11;
        weight_rom[609] = -32;
        weight_rom[610] = -28;
        weight_rom[611] = -28;
        weight_rom[612] = -14;
        weight_rom[613] = -14;
        weight_rom[614] = -11;
        weight_rom[615] = -2;
        weight_rom[616] = -2;
        weight_rom[617] = -2;
        weight_rom[618] = -13;
        weight_rom[619] = -12;
        weight_rom[620] = 20;
        weight_rom[621] = 23;
        weight_rom[622] = -6;
        weight_rom[623] = 12;
        weight_rom[624] = -8;
        weight_rom[625] = -9;
        weight_rom[626] = -6;
        weight_rom[627] = -6;
        weight_rom[628] = -6;
        weight_rom[629] = -13;
        weight_rom[630] = 0;
        weight_rom[631] = 1;
        weight_rom[632] = 3;
        weight_rom[633] = 5;
        weight_rom[634] = -14;
        weight_rom[635] = -18;
        weight_rom[636] = -20;
        weight_rom[637] = -40;
        weight_rom[638] = -31;
        weight_rom[639] = -36;
        weight_rom[640] = -20;
        weight_rom[641] = -28;
        weight_rom[642] = -4;
        weight_rom[643] = 2;
        weight_rom[644] = -1;
        weight_rom[645] = -3;
        weight_rom[646] = -12;
        weight_rom[647] = -26;
        weight_rom[648] = 28;
        weight_rom[649] = 24;
        weight_rom[650] = 15;
        weight_rom[651] = 7;
        weight_rom[652] = -14;
        weight_rom[653] = -2;
        weight_rom[654] = -4;
        weight_rom[655] = -4;
        weight_rom[656] = -10;
        weight_rom[657] = -10;
        weight_rom[658] = -4;
        weight_rom[659] = 0;
        weight_rom[660] = 2;
        weight_rom[661] = -9;
        weight_rom[662] = -23;
        weight_rom[663] = -23;
        weight_rom[664] = -25;
        weight_rom[665] = -38;
        weight_rom[666] = -23;
        weight_rom[667] = -28;
        weight_rom[668] = -15;
        weight_rom[669] = -25;
        weight_rom[670] = 14;
        weight_rom[671] = -4;
        weight_rom[672] = -3;
        weight_rom[673] = -4;
        weight_rom[674] = -7;
        weight_rom[675] = 20;
        weight_rom[676] = 5;
        weight_rom[677] = 24;
        weight_rom[678] = 15;
        weight_rom[679] = 16;
        weight_rom[680] = 15;
        weight_rom[681] = 9;
        weight_rom[682] = 0;
        weight_rom[683] = 8;
        weight_rom[684] = 1;
        weight_rom[685] = 8;
        weight_rom[686] = 1;
        weight_rom[687] = 3;
        weight_rom[688] = -10;
        weight_rom[689] = 1;
        weight_rom[690] = -6;
        weight_rom[691] = 1;
        weight_rom[692] = -5;
        weight_rom[693] = -15;
        weight_rom[694] = -34;
        weight_rom[695] = 0;
        weight_rom[696] = -15;
        weight_rom[697] = -25;
        weight_rom[698] = -3;
        weight_rom[699] = 3;
        weight_rom[700] = 4;
        weight_rom[701] = -1;
        weight_rom[702] = 4;
        weight_rom[703] = 15;
        weight_rom[704] = 15;
        weight_rom[705] = 5;
        weight_rom[706] = 12;
        weight_rom[707] = 15;
        weight_rom[708] = 37;
        weight_rom[709] = 32;
        weight_rom[710] = 25;
        weight_rom[711] = 34;
        weight_rom[712] = 47;
        weight_rom[713] = 21;
        weight_rom[714] = 20;
        weight_rom[715] = 24;
        weight_rom[716] = 29;
        weight_rom[717] = 32;
        weight_rom[718] = 32;
        weight_rom[719] = 17;
        weight_rom[720] = 8;
        weight_rom[721] = 9;
        weight_rom[722] = -1;
        weight_rom[723] = 7;
        weight_rom[724] = 10;
        weight_rom[725] = -4;
        weight_rom[726] = -3;
        weight_rom[727] = -4;
        weight_rom[728] = 2;
        weight_rom[729] = 4;
        weight_rom[730] = 3;
        weight_rom[731] = 2;
        weight_rom[732] = -18;
        weight_rom[733] = -11;
        weight_rom[734] = -10;
        weight_rom[735] = -2;
        weight_rom[736] = 8;
        weight_rom[737] = 27;
        weight_rom[738] = 20;
        weight_rom[739] = 31;
        weight_rom[740] = 16;
        weight_rom[741] = 41;
        weight_rom[742] = 36;
        weight_rom[743] = 39;
        weight_rom[744] = 29;
        weight_rom[745] = 44;
        weight_rom[746] = 25;
        weight_rom[747] = 31;
        weight_rom[748] = 14;
        weight_rom[749] = 0;
        weight_rom[750] = 25;
        weight_rom[751] = -4;
        weight_rom[752] = 1;
        weight_rom[753] = -1;
        weight_rom[754] = -4;
        weight_rom[755] = 1;
        weight_rom[756] = 3;
        weight_rom[757] = -4;
        weight_rom[758] = -2;
        weight_rom[759] = 3;
        weight_rom[760] = 0;
        weight_rom[761] = 17;
        weight_rom[762] = 20;
        weight_rom[763] = 25;
        weight_rom[764] = 24;
        weight_rom[765] = 6;
        weight_rom[766] = 27;
        weight_rom[767] = 7;
        weight_rom[768] = 18;
        weight_rom[769] = 32;
        weight_rom[770] = 21;
        weight_rom[771] = 7;
        weight_rom[772] = 18;
        weight_rom[773] = 29;
        weight_rom[774] = 16;
        weight_rom[775] = 7;
        weight_rom[776] = 3;
        weight_rom[777] = -16;
        weight_rom[778] = -3;
        weight_rom[779] = 3;
        weight_rom[780] = 3;
        weight_rom[781] = -4;
        weight_rom[782] = 1;
        weight_rom[783] = -2;
        weight_rom[784] = -4;
        weight_rom[785] = -4;
        weight_rom[786] = -1;
        weight_rom[787] = 4;
        weight_rom[788] = -4;
        weight_rom[789] = 4;
        weight_rom[790] = 4;
        weight_rom[791] = 3;
        weight_rom[792] = 4;
        weight_rom[793] = -1;
        weight_rom[794] = 4;
        weight_rom[795] = -3;
        weight_rom[796] = -4;
        weight_rom[797] = 12;
        weight_rom[798] = 1;
        weight_rom[799] = 0;
        weight_rom[800] = -1;
        weight_rom[801] = -3;
        weight_rom[802] = 2;
        weight_rom[803] = -2;
        weight_rom[804] = 3;
        weight_rom[805] = 1;
        weight_rom[806] = 4;
        weight_rom[807] = 0;
        weight_rom[808] = 2;
        weight_rom[809] = -2;
        weight_rom[810] = 1;
        weight_rom[811] = 3;
        weight_rom[812] = 2;
        weight_rom[813] = 1;
        weight_rom[814] = 1;
        weight_rom[815] = 3;
        weight_rom[816] = -1;
        weight_rom[817] = -1;
        weight_rom[818] = 16;
        weight_rom[819] = 24;
        weight_rom[820] = 15;
        weight_rom[821] = 21;
        weight_rom[822] = 26;
        weight_rom[823] = 34;
        weight_rom[824] = 43;
        weight_rom[825] = 36;
        weight_rom[826] = -2;
        weight_rom[827] = 11;
        weight_rom[828] = 1;
        weight_rom[829] = 16;
        weight_rom[830] = 27;
        weight_rom[831] = 22;
        weight_rom[832] = 23;
        weight_rom[833] = 16;
        weight_rom[834] = 20;
        weight_rom[835] = 15;
        weight_rom[836] = 0;
        weight_rom[837] = -1;
        weight_rom[838] = 2;
        weight_rom[839] = -1;
        weight_rom[840] = 3;
        weight_rom[841] = -3;
        weight_rom[842] = 1;
        weight_rom[843] = 1;
        weight_rom[844] = 12;
        weight_rom[845] = 3;
        weight_rom[846] = 20;
        weight_rom[847] = 42;
        weight_rom[848] = 43;
        weight_rom[849] = 24;
        weight_rom[850] = 50;
        weight_rom[851] = 29;
        weight_rom[852] = 41;
        weight_rom[853] = 24;
        weight_rom[854] = 21;
        weight_rom[855] = 19;
        weight_rom[856] = 2;
        weight_rom[857] = 17;
        weight_rom[858] = 23;
        weight_rom[859] = 18;
        weight_rom[860] = 22;
        weight_rom[861] = 10;
        weight_rom[862] = 32;
        weight_rom[863] = 22;
        weight_rom[864] = -4;
        weight_rom[865] = -14;
        weight_rom[866] = 4;
        weight_rom[867] = -3;
        weight_rom[868] = 3;
        weight_rom[869] = 2;
        weight_rom[870] = 11;
        weight_rom[871] = 4;
        weight_rom[872] = -2;
        weight_rom[873] = -14;
        weight_rom[874] = 13;
        weight_rom[875] = 3;
        weight_rom[876] = 1;
        weight_rom[877] = 24;
        weight_rom[878] = 5;
        weight_rom[879] = 4;
        weight_rom[880] = -2;
        weight_rom[881] = 3;
        weight_rom[882] = -11;
        weight_rom[883] = -7;
        weight_rom[884] = -9;
        weight_rom[885] = -8;
        weight_rom[886] = -5;
        weight_rom[887] = -11;
        weight_rom[888] = -5;
        weight_rom[889] = 24;
        weight_rom[890] = 30;
        weight_rom[891] = 26;
        weight_rom[892] = 20;
        weight_rom[893] = -30;
        weight_rom[894] = 0;
        weight_rom[895] = 0;
        weight_rom[896] = 1;
        weight_rom[897] = -4;
        weight_rom[898] = -11;
        weight_rom[899] = -2;
        weight_rom[900] = 8;
        weight_rom[901] = -21;
        weight_rom[902] = -22;
        weight_rom[903] = -6;
        weight_rom[904] = -12;
        weight_rom[905] = -4;
        weight_rom[906] = -5;
        weight_rom[907] = -7;
        weight_rom[908] = -7;
        weight_rom[909] = -3;
        weight_rom[910] = 3;
        weight_rom[911] = 1;
        weight_rom[912] = -8;
        weight_rom[913] = -1;
        weight_rom[914] = -17;
        weight_rom[915] = -6;
        weight_rom[916] = -11;
        weight_rom[917] = 9;
        weight_rom[918] = 4;
        weight_rom[919] = 25;
        weight_rom[920] = -9;
        weight_rom[921] = -7;
        weight_rom[922] = -11;
        weight_rom[923] = -2;
        weight_rom[924] = -4;
        weight_rom[925] = 1;
        weight_rom[926] = -4;
        weight_rom[927] = -18;
        weight_rom[928] = -17;
        weight_rom[929] = -45;
        weight_rom[930] = -33;
        weight_rom[931] = -24;
        weight_rom[932] = 1;
        weight_rom[933] = -10;
        weight_rom[934] = 4;
        weight_rom[935] = 9;
        weight_rom[936] = 6;
        weight_rom[937] = 18;
        weight_rom[938] = 19;
        weight_rom[939] = 10;
        weight_rom[940] = -5;
        weight_rom[941] = 5;
        weight_rom[942] = -2;
        weight_rom[943] = -2;
        weight_rom[944] = 1;
        weight_rom[945] = 13;
        weight_rom[946] = 0;
        weight_rom[947] = -4;
        weight_rom[948] = 23;
        weight_rom[949] = 12;
        weight_rom[950] = 15;
        weight_rom[951] = -3;
        weight_rom[952] = -4;
        weight_rom[953] = 4;
        weight_rom[954] = -2;
        weight_rom[955] = -35;
        weight_rom[956] = -32;
        weight_rom[957] = -33;
        weight_rom[958] = -36;
        weight_rom[959] = -5;
        weight_rom[960] = -2;
        weight_rom[961] = -11;
        weight_rom[962] = 2;
        weight_rom[963] = 9;
        weight_rom[964] = 16;
        weight_rom[965] = 13;
        weight_rom[966] = 21;
        weight_rom[967] = 24;
        weight_rom[968] = 16;
        weight_rom[969] = 17;
        weight_rom[970] = -4;
        weight_rom[971] = 0;
        weight_rom[972] = 4;
        weight_rom[973] = 2;
        weight_rom[974] = 8;
        weight_rom[975] = 9;
        weight_rom[976] = 10;
        weight_rom[977] = 18;
        weight_rom[978] = -7;
        weight_rom[979] = 14;
        weight_rom[980] = 3;
        weight_rom[981] = -17;
        weight_rom[982] = -1;
        weight_rom[983] = -44;
        weight_rom[984] = -32;
        weight_rom[985] = -39;
        weight_rom[986] = -29;
        weight_rom[987] = -13;
        weight_rom[988] = -3;
        weight_rom[989] = 4;
        weight_rom[990] = 1;
        weight_rom[991] = 14;
        weight_rom[992] = 16;
        weight_rom[993] = 10;
        weight_rom[994] = 13;
        weight_rom[995] = 32;
        weight_rom[996] = 19;
        weight_rom[997] = 6;
        weight_rom[998] = -2;
        weight_rom[999] = -13;
        weight_rom[1000] = -3;
        weight_rom[1001] = 7;
        weight_rom[1002] = 7;
        weight_rom[1003] = 16;
        weight_rom[1004] = 44;
        weight_rom[1005] = 10;
        weight_rom[1006] = -15;
        weight_rom[1007] = -4;
        weight_rom[1008] = 1;
        weight_rom[1009] = -16;
        weight_rom[1010] = -10;
        weight_rom[1011] = -41;
        weight_rom[1012] = -45;
        weight_rom[1013] = -30;
        weight_rom[1014] = -21;
        weight_rom[1015] = -16;
        weight_rom[1016] = 2;
        weight_rom[1017] = 3;
        weight_rom[1018] = 2;
        weight_rom[1019] = 7;
        weight_rom[1020] = 6;
        weight_rom[1021] = 10;
        weight_rom[1022] = 15;
        weight_rom[1023] = 14;
        weight_rom[1024] = 4;
        weight_rom[1025] = -31;
        weight_rom[1026] = -34;
        weight_rom[1027] = -16;
        weight_rom[1028] = -18;
        weight_rom[1029] = 9;
        weight_rom[1030] = -5;
        weight_rom[1031] = 22;
        weight_rom[1032] = 61;
        weight_rom[1033] = 2;
        weight_rom[1034] = -2;
        weight_rom[1035] = 16;
        weight_rom[1036] = -12;
        weight_rom[1037] = -25;
        weight_rom[1038] = -27;
        weight_rom[1039] = -37;
        weight_rom[1040] = -37;
        weight_rom[1041] = -18;
        weight_rom[1042] = -1;
        weight_rom[1043] = -2;
        weight_rom[1044] = 11;
        weight_rom[1045] = 10;
        weight_rom[1046] = 16;
        weight_rom[1047] = 23;
        weight_rom[1048] = 20;
        weight_rom[1049] = 23;
        weight_rom[1050] = 16;
        weight_rom[1051] = -12;
        weight_rom[1052] = -21;
        weight_rom[1053] = -42;
        weight_rom[1054] = -34;
        weight_rom[1055] = -18;
        weight_rom[1056] = -7;
        weight_rom[1057] = -2;
        weight_rom[1058] = -13;
        weight_rom[1059] = 23;
        weight_rom[1060] = 55;
        weight_rom[1061] = 0;
        weight_rom[1062] = -10;
        weight_rom[1063] = -16;
        weight_rom[1064] = -10;
        weight_rom[1065] = -14;
        weight_rom[1066] = -15;
        weight_rom[1067] = -57;
        weight_rom[1068] = -10;
        weight_rom[1069] = -8;
        weight_rom[1070] = -2;
        weight_rom[1071] = 12;
        weight_rom[1072] = 26;
        weight_rom[1073] = 37;
        weight_rom[1074] = 41;
        weight_rom[1075] = 44;
        weight_rom[1076] = 40;
        weight_rom[1077] = 29;
        weight_rom[1078] = 12;
        weight_rom[1079] = -24;
        weight_rom[1080] = -48;
        weight_rom[1081] = -45;
        weight_rom[1082] = -29;
        weight_rom[1083] = -13;
        weight_rom[1084] = -4;
        weight_rom[1085] = 2;
        weight_rom[1086] = 14;
        weight_rom[1087] = 41;
        weight_rom[1088] = 47;
        weight_rom[1089] = -46;
        weight_rom[1090] = -25;
        weight_rom[1091] = -11;
        weight_rom[1092] = 7;
        weight_rom[1093] = -12;
        weight_rom[1094] = -43;
        weight_rom[1095] = -44;
        weight_rom[1096] = -19;
        weight_rom[1097] = 8;
        weight_rom[1098] = 24;
        weight_rom[1099] = 36;
        weight_rom[1100] = 43;
        weight_rom[1101] = 49;
        weight_rom[1102] = 40;
        weight_rom[1103] = 37;
        weight_rom[1104] = 27;
        weight_rom[1105] = 32;
        weight_rom[1106] = 8;
        weight_rom[1107] = -21;
        weight_rom[1108] = -19;
        weight_rom[1109] = -27;
        weight_rom[1110] = -16;
        weight_rom[1111] = -6;
        weight_rom[1112] = 19;
        weight_rom[1113] = 41;
        weight_rom[1114] = 28;
        weight_rom[1115] = 45;
        weight_rom[1116] = 51;
        weight_rom[1117] = -21;
        weight_rom[1118] = -17;
        weight_rom[1119] = 12;
        weight_rom[1120] = 7;
        weight_rom[1121] = -14;
        weight_rom[1122] = -24;
        weight_rom[1123] = -23;
        weight_rom[1124] = 7;
        weight_rom[1125] = 33;
        weight_rom[1126] = 50;
        weight_rom[1127] = 39;
        weight_rom[1128] = 44;
        weight_rom[1129] = 45;
        weight_rom[1130] = 29;
        weight_rom[1131] = 30;
        weight_rom[1132] = 10;
        weight_rom[1133] = 24;
        weight_rom[1134] = 5;
        weight_rom[1135] = -9;
        weight_rom[1136] = -14;
        weight_rom[1137] = -4;
        weight_rom[1138] = -9;
        weight_rom[1139] = 14;
        weight_rom[1140] = 22;
        weight_rom[1141] = 52;
        weight_rom[1142] = 63;
        weight_rom[1143] = 65;
        weight_rom[1144] = 50;
        weight_rom[1145] = -29;
        weight_rom[1146] = -49;
        weight_rom[1147] = 14;
        weight_rom[1148] = 4;
        weight_rom[1149] = -10;
        weight_rom[1150] = -27;
        weight_rom[1151] = 7;
        weight_rom[1152] = 6;
        weight_rom[1153] = 45;
        weight_rom[1154] = 52;
        weight_rom[1155] = 47;
        weight_rom[1156] = 33;
        weight_rom[1157] = 33;
        weight_rom[1158] = 27;
        weight_rom[1159] = 16;
        weight_rom[1160] = 12;
        weight_rom[1161] = 0;
        weight_rom[1162] = 2;
        weight_rom[1163] = 10;
        weight_rom[1164] = 2;
        weight_rom[1165] = -9;
        weight_rom[1166] = -5;
        weight_rom[1167] = 13;
        weight_rom[1168] = 28;
        weight_rom[1169] = 39;
        weight_rom[1170] = 56;
        weight_rom[1171] = 64;
        weight_rom[1172] = 26;
        weight_rom[1173] = -21;
        weight_rom[1174] = -54;
        weight_rom[1175] = -25;
        weight_rom[1176] = 0;
        weight_rom[1177] = -2;
        weight_rom[1178] = -18;
        weight_rom[1179] = -3;
        weight_rom[1180] = 11;
        weight_rom[1181] = 36;
        weight_rom[1182] = 35;
        weight_rom[1183] = 37;
        weight_rom[1184] = 19;
        weight_rom[1185] = 14;
        weight_rom[1186] = 23;
        weight_rom[1187] = 26;
        weight_rom[1188] = 0;
        weight_rom[1189] = 10;
        weight_rom[1190] = 0;
        weight_rom[1191] = 7;
        weight_rom[1192] = 7;
        weight_rom[1193] = -7;
        weight_rom[1194] = -6;
        weight_rom[1195] = -5;
        weight_rom[1196] = 2;
        weight_rom[1197] = 23;
        weight_rom[1198] = 31;
        weight_rom[1199] = 24;
        weight_rom[1200] = 20;
        weight_rom[1201] = -17;
        weight_rom[1202] = -32;
        weight_rom[1203] = 2;
        weight_rom[1204] = -3;
        weight_rom[1205] = -13;
        weight_rom[1206] = -28;
        weight_rom[1207] = -12;
        weight_rom[1208] = -19;
        weight_rom[1209] = 10;
        weight_rom[1210] = 5;
        weight_rom[1211] = 20;
        weight_rom[1212] = 15;
        weight_rom[1213] = 16;
        weight_rom[1214] = 18;
        weight_rom[1215] = 14;
        weight_rom[1216] = 2;
        weight_rom[1217] = -2;
        weight_rom[1218] = -1;
        weight_rom[1219] = -8;
        weight_rom[1220] = -2;
        weight_rom[1221] = -6;
        weight_rom[1222] = -2;
        weight_rom[1223] = -14;
        weight_rom[1224] = 9;
        weight_rom[1225] = 7;
        weight_rom[1226] = -1;
        weight_rom[1227] = 7;
        weight_rom[1228] = 4;
        weight_rom[1229] = -2;
        weight_rom[1230] = -40;
        weight_rom[1231] = -17;
        weight_rom[1232] = 3;
        weight_rom[1233] = -1;
        weight_rom[1234] = -22;
        weight_rom[1235] = -24;
        weight_rom[1236] = -37;
        weight_rom[1237] = -9;
        weight_rom[1238] = 5;
        weight_rom[1239] = 10;
        weight_rom[1240] = 16;
        weight_rom[1241] = 4;
        weight_rom[1242] = 20;
        weight_rom[1243] = 22;
        weight_rom[1244] = -1;
        weight_rom[1245] = -24;
        weight_rom[1246] = -13;
        weight_rom[1247] = -8;
        weight_rom[1248] = 1;
        weight_rom[1249] = -10;
        weight_rom[1250] = -11;
        weight_rom[1251] = -16;
        weight_rom[1252] = -3;
        weight_rom[1253] = -6;
        weight_rom[1254] = -4;
        weight_rom[1255] = -8;
        weight_rom[1256] = -17;
        weight_rom[1257] = -25;
        weight_rom[1258] = -51;
        weight_rom[1259] = -22;
        weight_rom[1260] = -2;
        weight_rom[1261] = 2;
        weight_rom[1262] = -29;
        weight_rom[1263] = -35;
        weight_rom[1264] = -61;
        weight_rom[1265] = -17;
        weight_rom[1266] = -7;
        weight_rom[1267] = -1;
        weight_rom[1268] = 11;
        weight_rom[1269] = 25;
        weight_rom[1270] = 35;
        weight_rom[1271] = 23;
        weight_rom[1272] = 2;
        weight_rom[1273] = -10;
        weight_rom[1274] = -5;
        weight_rom[1275] = -1;
        weight_rom[1276] = 6;
        weight_rom[1277] = -2;
        weight_rom[1278] = -5;
        weight_rom[1279] = -4;
        weight_rom[1280] = -1;
        weight_rom[1281] = -6;
        weight_rom[1282] = 0;
        weight_rom[1283] = -14;
        weight_rom[1284] = 14;
        weight_rom[1285] = -17;
        weight_rom[1286] = -39;
        weight_rom[1287] = 4;
        weight_rom[1288] = 0;
        weight_rom[1289] = -1;
        weight_rom[1290] = -18;
        weight_rom[1291] = -40;
        weight_rom[1292] = -46;
        weight_rom[1293] = -42;
        weight_rom[1294] = -22;
        weight_rom[1295] = 11;
        weight_rom[1296] = 17;
        weight_rom[1297] = 22;
        weight_rom[1298] = 31;
        weight_rom[1299] = 22;
        weight_rom[1300] = 12;
        weight_rom[1301] = 2;
        weight_rom[1302] = -2;
        weight_rom[1303] = 2;
        weight_rom[1304] = -2;
        weight_rom[1305] = -6;
        weight_rom[1306] = 6;
        weight_rom[1307] = -3;
        weight_rom[1308] = 6;
        weight_rom[1309] = -3;
        weight_rom[1310] = -2;
        weight_rom[1311] = 3;
        weight_rom[1312] = -5;
        weight_rom[1313] = -9;
        weight_rom[1314] = -10;
        weight_rom[1315] = -19;
        weight_rom[1316] = 2;
        weight_rom[1317] = 1;
        weight_rom[1318] = 2;
        weight_rom[1319] = -44;
        weight_rom[1320] = -34;
        weight_rom[1321] = -24;
        weight_rom[1322] = -4;
        weight_rom[1323] = 7;
        weight_rom[1324] = -1;
        weight_rom[1325] = 13;
        weight_rom[1326] = 27;
        weight_rom[1327] = 21;
        weight_rom[1328] = 16;
        weight_rom[1329] = 2;
        weight_rom[1330] = 5;
        weight_rom[1331] = 5;
        weight_rom[1332] = -2;
        weight_rom[1333] = -8;
        weight_rom[1334] = -1;
        weight_rom[1335] = 5;
        weight_rom[1336] = 20;
        weight_rom[1337] = 3;
        weight_rom[1338] = 12;
        weight_rom[1339] = 9;
        weight_rom[1340] = -4;
        weight_rom[1341] = -31;
        weight_rom[1342] = -25;
        weight_rom[1343] = -5;
        weight_rom[1344] = -3;
        weight_rom[1345] = 10;
        weight_rom[1346] = -8;
        weight_rom[1347] = -25;
        weight_rom[1348] = -16;
        weight_rom[1349] = -5;
        weight_rom[1350] = -13;
        weight_rom[1351] = -4;
        weight_rom[1352] = 7;
        weight_rom[1353] = 7;
        weight_rom[1354] = 19;
        weight_rom[1355] = 16;
        weight_rom[1356] = 20;
        weight_rom[1357] = 22;
        weight_rom[1358] = 15;
        weight_rom[1359] = 10;
        weight_rom[1360] = 4;
        weight_rom[1361] = -4;
        weight_rom[1362] = 10;
        weight_rom[1363] = 8;
        weight_rom[1364] = 1;
        weight_rom[1365] = 2;
        weight_rom[1366] = 8;
        weight_rom[1367] = 3;
        weight_rom[1368] = -34;
        weight_rom[1369] = -15;
        weight_rom[1370] = -6;
        weight_rom[1371] = -4;
        weight_rom[1372] = -3;
        weight_rom[1373] = 2;
        weight_rom[1374] = -2;
        weight_rom[1375] = -30;
        weight_rom[1376] = -11;
        weight_rom[1377] = 4;
        weight_rom[1378] = 3;
        weight_rom[1379] = 3;
        weight_rom[1380] = 5;
        weight_rom[1381] = 19;
        weight_rom[1382] = 19;
        weight_rom[1383] = 18;
        weight_rom[1384] = 30;
        weight_rom[1385] = 27;
        weight_rom[1386] = 26;
        weight_rom[1387] = 22;
        weight_rom[1388] = 8;
        weight_rom[1389] = 7;
        weight_rom[1390] = 2;
        weight_rom[1391] = -10;
        weight_rom[1392] = 5;
        weight_rom[1393] = -2;
        weight_rom[1394] = 4;
        weight_rom[1395] = -7;
        weight_rom[1396] = -17;
        weight_rom[1397] = -11;
        weight_rom[1398] = 6;
        weight_rom[1399] = 4;
        weight_rom[1400] = -1;
        weight_rom[1401] = -3;
        weight_rom[1402] = -15;
        weight_rom[1403] = -35;
        weight_rom[1404] = -10;
        weight_rom[1405] = -12;
        weight_rom[1406] = -2;
        weight_rom[1407] = 5;
        weight_rom[1408] = 9;
        weight_rom[1409] = 6;
        weight_rom[1410] = 25;
        weight_rom[1411] = 15;
        weight_rom[1412] = 27;
        weight_rom[1413] = 33;
        weight_rom[1414] = 33;
        weight_rom[1415] = 19;
        weight_rom[1416] = 14;
        weight_rom[1417] = -2;
        weight_rom[1418] = 1;
        weight_rom[1419] = -11;
        weight_rom[1420] = -4;
        weight_rom[1421] = -6;
        weight_rom[1422] = -6;
        weight_rom[1423] = 3;
        weight_rom[1424] = -2;
        weight_rom[1425] = -6;
        weight_rom[1426] = -1;
        weight_rom[1427] = -2;
        weight_rom[1428] = 1;
        weight_rom[1429] = -3;
        weight_rom[1430] = -23;
        weight_rom[1431] = -21;
        weight_rom[1432] = -30;
        weight_rom[1433] = -14;
        weight_rom[1434] = -22;
        weight_rom[1435] = -17;
        weight_rom[1436] = 9;
        weight_rom[1437] = 0;
        weight_rom[1438] = 9;
        weight_rom[1439] = 8;
        weight_rom[1440] = 26;
        weight_rom[1441] = 24;
        weight_rom[1442] = 27;
        weight_rom[1443] = 14;
        weight_rom[1444] = 16;
        weight_rom[1445] = 6;
        weight_rom[1446] = -4;
        weight_rom[1447] = -4;
        weight_rom[1448] = -7;
        weight_rom[1449] = 5;
        weight_rom[1450] = 7;
        weight_rom[1451] = 23;
        weight_rom[1452] = 11;
        weight_rom[1453] = -8;
        weight_rom[1454] = -8;
        weight_rom[1455] = 3;
        weight_rom[1456] = -4;
        weight_rom[1457] = 0;
        weight_rom[1458] = -6;
        weight_rom[1459] = -33;
        weight_rom[1460] = -46;
        weight_rom[1461] = -30;
        weight_rom[1462] = -30;
        weight_rom[1463] = -33;
        weight_rom[1464] = -11;
        weight_rom[1465] = -4;
        weight_rom[1466] = 4;
        weight_rom[1467] = -8;
        weight_rom[1468] = 8;
        weight_rom[1469] = -7;
        weight_rom[1470] = 0;
        weight_rom[1471] = 11;
        weight_rom[1472] = 4;
        weight_rom[1473] = -8;
        weight_rom[1474] = 11;
        weight_rom[1475] = 11;
        weight_rom[1476] = 15;
        weight_rom[1477] = -7;
        weight_rom[1478] = 10;
        weight_rom[1479] = 27;
        weight_rom[1480] = 7;
        weight_rom[1481] = -5;
        weight_rom[1482] = -3;
        weight_rom[1483] = -1;
        weight_rom[1484] = 0;
        weight_rom[1485] = -1;
        weight_rom[1486] = -3;
        weight_rom[1487] = 4;
        weight_rom[1488] = -20;
        weight_rom[1489] = -30;
        weight_rom[1490] = -38;
        weight_rom[1491] = -28;
        weight_rom[1492] = -52;
        weight_rom[1493] = -36;
        weight_rom[1494] = -31;
        weight_rom[1495] = -28;
        weight_rom[1496] = -25;
        weight_rom[1497] = -19;
        weight_rom[1498] = -16;
        weight_rom[1499] = -7;
        weight_rom[1500] = 0;
        weight_rom[1501] = 0;
        weight_rom[1502] = 11;
        weight_rom[1503] = 13;
        weight_rom[1504] = 36;
        weight_rom[1505] = 22;
        weight_rom[1506] = 3;
        weight_rom[1507] = 22;
        weight_rom[1508] = 12;
        weight_rom[1509] = 4;
        weight_rom[1510] = 1;
        weight_rom[1511] = 3;
        weight_rom[1512] = 3;
        weight_rom[1513] = 0;
        weight_rom[1514] = 1;
        weight_rom[1515] = 0;
        weight_rom[1516] = 25;
        weight_rom[1517] = 19;
        weight_rom[1518] = 6;
        weight_rom[1519] = -8;
        weight_rom[1520] = -6;
        weight_rom[1521] = -7;
        weight_rom[1522] = -5;
        weight_rom[1523] = 3;
        weight_rom[1524] = 12;
        weight_rom[1525] = 1;
        weight_rom[1526] = 16;
        weight_rom[1527] = -5;
        weight_rom[1528] = -1;
        weight_rom[1529] = -5;
        weight_rom[1530] = 10;
        weight_rom[1531] = -2;
        weight_rom[1532] = 15;
        weight_rom[1533] = 22;
        weight_rom[1534] = -6;
        weight_rom[1535] = 9;
        weight_rom[1536] = 2;
        weight_rom[1537] = 0;
        weight_rom[1538] = 3;
        weight_rom[1539] = 1;
        weight_rom[1540] = -3;
        weight_rom[1541] = 1;
        weight_rom[1542] = 3;
        weight_rom[1543] = -3;
        weight_rom[1544] = 4;
        weight_rom[1545] = -24;
        weight_rom[1546] = -24;
        weight_rom[1547] = 7;
        weight_rom[1548] = 5;
        weight_rom[1549] = -3;
        weight_rom[1550] = -11;
        weight_rom[1551] = 3;
        weight_rom[1552] = -2;
        weight_rom[1553] = -34;
        weight_rom[1554] = -5;
        weight_rom[1555] = 0;
        weight_rom[1556] = -1;
        weight_rom[1557] = -28;
        weight_rom[1558] = -4;
        weight_rom[1559] = 10;
        weight_rom[1560] = -4;
        weight_rom[1561] = -3;
        weight_rom[1562] = -6;
        weight_rom[1563] = 3;
        weight_rom[1564] = 4;
        weight_rom[1565] = -4;
        weight_rom[1566] = 1;
        weight_rom[1567] = -4;
        weight_rom[1568] = -3;
        weight_rom[1569] = 3;
        weight_rom[1570] = 4;
        weight_rom[1571] = 3;
        weight_rom[1572] = 1;
        weight_rom[1573] = -2;
        weight_rom[1574] = 4;
        weight_rom[1575] = -2;
        weight_rom[1576] = -1;
        weight_rom[1577] = 1;
        weight_rom[1578] = 3;
        weight_rom[1579] = 3;
        weight_rom[1580] = 4;
        weight_rom[1581] = -12;
        weight_rom[1582] = -8;
        weight_rom[1583] = 3;
        weight_rom[1584] = 4;
        weight_rom[1585] = 4;
        weight_rom[1586] = -2;
        weight_rom[1587] = 3;
        weight_rom[1588] = -2;
        weight_rom[1589] = 4;
        weight_rom[1590] = -4;
        weight_rom[1591] = 2;
        weight_rom[1592] = -2;
        weight_rom[1593] = -4;
        weight_rom[1594] = -3;
        weight_rom[1595] = -4;
        weight_rom[1596] = -5;
        weight_rom[1597] = 1;
        weight_rom[1598] = 1;
        weight_rom[1599] = 0;
        weight_rom[1600] = -4;
        weight_rom[1601] = -1;
        weight_rom[1602] = -14;
        weight_rom[1603] = -24;
        weight_rom[1604] = -24;
        weight_rom[1605] = -24;
        weight_rom[1606] = -25;
        weight_rom[1607] = -26;
        weight_rom[1608] = -36;
        weight_rom[1609] = -28;
        weight_rom[1610] = -1;
        weight_rom[1611] = -25;
        weight_rom[1612] = -32;
        weight_rom[1613] = -32;
        weight_rom[1614] = -26;
        weight_rom[1615] = -20;
        weight_rom[1616] = -18;
        weight_rom[1617] = -18;
        weight_rom[1618] = -19;
        weight_rom[1619] = -14;
        weight_rom[1620] = 2;
        weight_rom[1621] = -3;
        weight_rom[1622] = 1;
        weight_rom[1623] = 3;
        weight_rom[1624] = 4;
        weight_rom[1625] = 3;
        weight_rom[1626] = 0;
        weight_rom[1627] = 3;
        weight_rom[1628] = -13;
        weight_rom[1629] = -4;
        weight_rom[1630] = -22;
        weight_rom[1631] = -43;
        weight_rom[1632] = -33;
        weight_rom[1633] = -42;
        weight_rom[1634] = -52;
        weight_rom[1635] = -59;
        weight_rom[1636] = -71;
        weight_rom[1637] = -50;
        weight_rom[1638] = -45;
        weight_rom[1639] = -46;
        weight_rom[1640] = -38;
        weight_rom[1641] = -48;
        weight_rom[1642] = -23;
        weight_rom[1643] = -17;
        weight_rom[1644] = -27;
        weight_rom[1645] = -26;
        weight_rom[1646] = -18;
        weight_rom[1647] = -20;
        weight_rom[1648] = -16;
        weight_rom[1649] = -7;
        weight_rom[1650] = -3;
        weight_rom[1651] = 2;
        weight_rom[1652] = 1;
        weight_rom[1653] = -3;
        weight_rom[1654] = -9;
        weight_rom[1655] = -1;
        weight_rom[1656] = 4;
        weight_rom[1657] = 5;
        weight_rom[1658] = -35;
        weight_rom[1659] = -37;
        weight_rom[1660] = -41;
        weight_rom[1661] = -75;
        weight_rom[1662] = -36;
        weight_rom[1663] = -45;
        weight_rom[1664] = -60;
        weight_rom[1665] = -61;
        weight_rom[1666] = -37;
        weight_rom[1667] = -36;
        weight_rom[1668] = -27;
        weight_rom[1669] = -23;
        weight_rom[1670] = -8;
        weight_rom[1671] = -14;
        weight_rom[1672] = -11;
        weight_rom[1673] = -10;
        weight_rom[1674] = -26;
        weight_rom[1675] = -10;
        weight_rom[1676] = -12;
        weight_rom[1677] = -9;
        weight_rom[1678] = 3;
        weight_rom[1679] = -1;
        weight_rom[1680] = -1;
        weight_rom[1681] = 1;
        weight_rom[1682] = -8;
        weight_rom[1683] = -4;
        weight_rom[1684] = 4;
        weight_rom[1685] = 6;
        weight_rom[1686] = -6;
        weight_rom[1687] = -8;
        weight_rom[1688] = -16;
        weight_rom[1689] = -16;
        weight_rom[1690] = -15;
        weight_rom[1691] = -9;
        weight_rom[1692] = -4;
        weight_rom[1693] = -9;
        weight_rom[1694] = -4;
        weight_rom[1695] = 0;
        weight_rom[1696] = 2;
        weight_rom[1697] = -14;
        weight_rom[1698] = -9;
        weight_rom[1699] = -2;
        weight_rom[1700] = 1;
        weight_rom[1701] = -11;
        weight_rom[1702] = -18;
        weight_rom[1703] = -8;
        weight_rom[1704] = 24;
        weight_rom[1705] = 27;
        weight_rom[1706] = 20;
        weight_rom[1707] = 4;
        weight_rom[1708] = 1;
        weight_rom[1709] = -1;
        weight_rom[1710] = -3;
        weight_rom[1711] = 0;
        weight_rom[1712] = -11;
        weight_rom[1713] = 5;
        weight_rom[1714] = -12;
        weight_rom[1715] = 1;
        weight_rom[1716] = -12;
        weight_rom[1717] = -7;
        weight_rom[1718] = -27;
        weight_rom[1719] = 9;
        weight_rom[1720] = 11;
        weight_rom[1721] = 5;
        weight_rom[1722] = 2;
        weight_rom[1723] = 4;
        weight_rom[1724] = 4;
        weight_rom[1725] = 0;
        weight_rom[1726] = -13;
        weight_rom[1727] = 1;
        weight_rom[1728] = -7;
        weight_rom[1729] = -27;
        weight_rom[1730] = -26;
        weight_rom[1731] = -21;
        weight_rom[1732] = -12;
        weight_rom[1733] = 9;
        weight_rom[1734] = 5;
        weight_rom[1735] = -1;
        weight_rom[1736] = -2;
        weight_rom[1737] = -4;
        weight_rom[1738] = 13;
        weight_rom[1739] = 2;
        weight_rom[1740] = 7;
        weight_rom[1741] = -6;
        weight_rom[1742] = 6;
        weight_rom[1743] = -10;
        weight_rom[1744] = 10;
        weight_rom[1745] = 6;
        weight_rom[1746] = 7;
        weight_rom[1747] = 13;
        weight_rom[1748] = 16;
        weight_rom[1749] = 22;
        weight_rom[1750] = 27;
        weight_rom[1751] = 32;
        weight_rom[1752] = 17;
        weight_rom[1753] = 23;
        weight_rom[1754] = 5;
        weight_rom[1755] = 9;
        weight_rom[1756] = 5;
        weight_rom[1757] = -4;
        weight_rom[1758] = -10;
        weight_rom[1759] = -3;
        weight_rom[1760] = -6;
        weight_rom[1761] = 20;
        weight_rom[1762] = -13;
        weight_rom[1763] = -5;
        weight_rom[1764] = 0;
        weight_rom[1765] = 4;
        weight_rom[1766] = -25;
        weight_rom[1767] = 11;
        weight_rom[1768] = -4;
        weight_rom[1769] = 0;
        weight_rom[1770] = -1;
        weight_rom[1771] = 1;
        weight_rom[1772] = 8;
        weight_rom[1773] = 8;
        weight_rom[1774] = 1;
        weight_rom[1775] = 3;
        weight_rom[1776] = 21;
        weight_rom[1777] = 26;
        weight_rom[1778] = 25;
        weight_rom[1779] = 36;
        weight_rom[1780] = 19;
        weight_rom[1781] = 25;
        weight_rom[1782] = 11;
        weight_rom[1783] = 12;
        weight_rom[1784] = 5;
        weight_rom[1785] = 5;
        weight_rom[1786] = -13;
        weight_rom[1787] = 6;
        weight_rom[1788] = 8;
        weight_rom[1789] = 7;
        weight_rom[1790] = -5;
        weight_rom[1791] = 4;
        weight_rom[1792] = -13;
        weight_rom[1793] = -12;
        weight_rom[1794] = 2;
        weight_rom[1795] = 0;
        weight_rom[1796] = 2;
        weight_rom[1797] = 3;
        weight_rom[1798] = 10;
        weight_rom[1799] = 5;
        weight_rom[1800] = 5;
        weight_rom[1801] = 7;
        weight_rom[1802] = -4;
        weight_rom[1803] = 6;
        weight_rom[1804] = 11;
        weight_rom[1805] = 20;
        weight_rom[1806] = 11;
        weight_rom[1807] = 9;
        weight_rom[1808] = 22;
        weight_rom[1809] = 5;
        weight_rom[1810] = 22;
        weight_rom[1811] = 1;
        weight_rom[1812] = 5;
        weight_rom[1813] = 13;
        weight_rom[1814] = 9;
        weight_rom[1815] = -3;
        weight_rom[1816] = 33;
        weight_rom[1817] = 21;
        weight_rom[1818] = 22;
        weight_rom[1819] = 11;
        weight_rom[1820] = -6;
        weight_rom[1821] = -7;
        weight_rom[1822] = -8;
        weight_rom[1823] = -2;
        weight_rom[1824] = 4;
        weight_rom[1825] = 3;
        weight_rom[1826] = 18;
        weight_rom[1827] = 15;
        weight_rom[1828] = 2;
        weight_rom[1829] = 11;
        weight_rom[1830] = -6;
        weight_rom[1831] = -4;
        weight_rom[1832] = 3;
        weight_rom[1833] = 4;
        weight_rom[1834] = -4;
        weight_rom[1835] = -6;
        weight_rom[1836] = 0;
        weight_rom[1837] = 8;
        weight_rom[1838] = 8;
        weight_rom[1839] = 17;
        weight_rom[1840] = 17;
        weight_rom[1841] = 19;
        weight_rom[1842] = 22;
        weight_rom[1843] = 13;
        weight_rom[1844] = -3;
        weight_rom[1845] = 12;
        weight_rom[1846] = 12;
        weight_rom[1847] = -11;
        weight_rom[1848] = -16;
        weight_rom[1849] = -23;
        weight_rom[1850] = -38;
        weight_rom[1851] = 14;
        weight_rom[1852] = 7;
        weight_rom[1853] = 3;
        weight_rom[1854] = 16;
        weight_rom[1855] = 14;
        weight_rom[1856] = 13;
        weight_rom[1857] = 6;
        weight_rom[1858] = -3;
        weight_rom[1859] = -6;
        weight_rom[1860] = -6;
        weight_rom[1861] = -14;
        weight_rom[1862] = -17;
        weight_rom[1863] = -18;
        weight_rom[1864] = 5;
        weight_rom[1865] = -3;
        weight_rom[1866] = 11;
        weight_rom[1867] = 24;
        weight_rom[1868] = 20;
        weight_rom[1869] = 20;
        weight_rom[1870] = 14;
        weight_rom[1871] = 8;
        weight_rom[1872] = -28;
        weight_rom[1873] = -20;
        weight_rom[1874] = -14;
        weight_rom[1875] = 8;
        weight_rom[1876] = -22;
        weight_rom[1877] = -11;
        weight_rom[1878] = -37;
        weight_rom[1879] = 26;
        weight_rom[1880] = 16;
        weight_rom[1881] = 18;
        weight_rom[1882] = 20;
        weight_rom[1883] = 9;
        weight_rom[1884] = 9;
        weight_rom[1885] = 15;
        weight_rom[1886] = 17;
        weight_rom[1887] = 19;
        weight_rom[1888] = 23;
        weight_rom[1889] = 0;
        weight_rom[1890] = 5;
        weight_rom[1891] = 18;
        weight_rom[1892] = 13;
        weight_rom[1893] = 22;
        weight_rom[1894] = 10;
        weight_rom[1895] = 15;
        weight_rom[1896] = 23;
        weight_rom[1897] = 16;
        weight_rom[1898] = 21;
        weight_rom[1899] = -9;
        weight_rom[1900] = -2;
        weight_rom[1901] = 0;
        weight_rom[1902] = 19;
        weight_rom[1903] = -1;
        weight_rom[1904] = -12;
        weight_rom[1905] = -11;
        weight_rom[1906] = -25;
        weight_rom[1907] = 13;
        weight_rom[1908] = 27;
        weight_rom[1909] = 25;
        weight_rom[1910] = 17;
        weight_rom[1911] = 25;
        weight_rom[1912] = 21;
        weight_rom[1913] = 23;
        weight_rom[1914] = 18;
        weight_rom[1915] = 25;
        weight_rom[1916] = 22;
        weight_rom[1917] = 20;
        weight_rom[1918] = 14;
        weight_rom[1919] = 22;
        weight_rom[1920] = 19;
        weight_rom[1921] = 26;
        weight_rom[1922] = 20;
        weight_rom[1923] = 24;
        weight_rom[1924] = 24;
        weight_rom[1925] = 19;
        weight_rom[1926] = 18;
        weight_rom[1927] = 3;
        weight_rom[1928] = -9;
        weight_rom[1929] = -5;
        weight_rom[1930] = -8;
        weight_rom[1931] = 4;
        weight_rom[1932] = 0;
        weight_rom[1933] = 0;
        weight_rom[1934] = -27;
        weight_rom[1935] = 13;
        weight_rom[1936] = 34;
        weight_rom[1937] = 30;
        weight_rom[1938] = 27;
        weight_rom[1939] = 41;
        weight_rom[1940] = 26;
        weight_rom[1941] = 29;
        weight_rom[1942] = 17;
        weight_rom[1943] = 20;
        weight_rom[1944] = 5;
        weight_rom[1945] = 18;
        weight_rom[1946] = 13;
        weight_rom[1947] = 29;
        weight_rom[1948] = 32;
        weight_rom[1949] = 22;
        weight_rom[1950] = 31;
        weight_rom[1951] = 23;
        weight_rom[1952] = 18;
        weight_rom[1953] = 13;
        weight_rom[1954] = -6;
        weight_rom[1955] = -22;
        weight_rom[1956] = -24;
        weight_rom[1957] = -15;
        weight_rom[1958] = -12;
        weight_rom[1959] = -15;
        weight_rom[1960] = 4;
        weight_rom[1961] = -5;
        weight_rom[1962] = -12;
        weight_rom[1963] = 20;
        weight_rom[1964] = 40;
        weight_rom[1965] = 8;
        weight_rom[1966] = 20;
        weight_rom[1967] = 7;
        weight_rom[1968] = 18;
        weight_rom[1969] = 5;
        weight_rom[1970] = 7;
        weight_rom[1971] = 4;
        weight_rom[1972] = 11;
        weight_rom[1973] = 13;
        weight_rom[1974] = 12;
        weight_rom[1975] = 16;
        weight_rom[1976] = 18;
        weight_rom[1977] = 35;
        weight_rom[1978] = 28;
        weight_rom[1979] = 24;
        weight_rom[1980] = 0;
        weight_rom[1981] = 0;
        weight_rom[1982] = -20;
        weight_rom[1983] = -36;
        weight_rom[1984] = -44;
        weight_rom[1985] = -26;
        weight_rom[1986] = -41;
        weight_rom[1987] = 3;
        weight_rom[1988] = 1;
        weight_rom[1989] = 5;
        weight_rom[1990] = 7;
        weight_rom[1991] = 11;
        weight_rom[1992] = 9;
        weight_rom[1993] = -14;
        weight_rom[1994] = 3;
        weight_rom[1995] = 5;
        weight_rom[1996] = 1;
        weight_rom[1997] = 3;
        weight_rom[1998] = 9;
        weight_rom[1999] = 1;
        weight_rom[2000] = 16;
        weight_rom[2001] = 14;
        weight_rom[2002] = 11;
        weight_rom[2003] = 21;
        weight_rom[2004] = 18;
        weight_rom[2005] = 31;
        weight_rom[2006] = 14;
        weight_rom[2007] = 12;
        weight_rom[2008] = 11;
        weight_rom[2009] = -4;
        weight_rom[2010] = 4;
        weight_rom[2011] = -18;
        weight_rom[2012] = -63;
        weight_rom[2013] = -42;
        weight_rom[2014] = -12;
        weight_rom[2015] = -13;
        weight_rom[2016] = -2;
        weight_rom[2017] = -3;
        weight_rom[2018] = 30;
        weight_rom[2019] = 0;
        weight_rom[2020] = -11;
        weight_rom[2021] = -27;
        weight_rom[2022] = 1;
        weight_rom[2023] = 9;
        weight_rom[2024] = 18;
        weight_rom[2025] = 9;
        weight_rom[2026] = 8;
        weight_rom[2027] = 8;
        weight_rom[2028] = 28;
        weight_rom[2029] = 11;
        weight_rom[2030] = 2;
        weight_rom[2031] = 8;
        weight_rom[2032] = 15;
        weight_rom[2033] = 21;
        weight_rom[2034] = 19;
        weight_rom[2035] = 2;
        weight_rom[2036] = -10;
        weight_rom[2037] = -24;
        weight_rom[2038] = -14;
        weight_rom[2039] = -1;
        weight_rom[2040] = -34;
        weight_rom[2041] = -58;
        weight_rom[2042] = -38;
        weight_rom[2043] = -6;
        weight_rom[2044] = -2;
        weight_rom[2045] = 9;
        weight_rom[2046] = 0;
        weight_rom[2047] = 6;
        weight_rom[2048] = -5;
        weight_rom[2049] = -14;
        weight_rom[2050] = -20;
        weight_rom[2051] = 2;
        weight_rom[2052] = 8;
        weight_rom[2053] = 8;
        weight_rom[2054] = -6;
        weight_rom[2055] = -3;
        weight_rom[2056] = 21;
        weight_rom[2057] = 9;
        weight_rom[2058] = -1;
        weight_rom[2059] = 7;
        weight_rom[2060] = 18;
        weight_rom[2061] = 16;
        weight_rom[2062] = 9;
        weight_rom[2063] = 6;
        weight_rom[2064] = -3;
        weight_rom[2065] = 10;
        weight_rom[2066] = -9;
        weight_rom[2067] = -5;
        weight_rom[2068] = -32;
        weight_rom[2069] = -63;
        weight_rom[2070] = -34;
        weight_rom[2071] = -2;
        weight_rom[2072] = -1;
        weight_rom[2073] = 5;
        weight_rom[2074] = 2;
        weight_rom[2075] = 10;
        weight_rom[2076] = -9;
        weight_rom[2077] = -13;
        weight_rom[2078] = -11;
        weight_rom[2079] = -15;
        weight_rom[2080] = -17;
        weight_rom[2081] = -13;
        weight_rom[2082] = -9;
        weight_rom[2083] = -9;
        weight_rom[2084] = -17;
        weight_rom[2085] = -14;
        weight_rom[2086] = -16;
        weight_rom[2087] = 4;
        weight_rom[2088] = 8;
        weight_rom[2089] = 4;
        weight_rom[2090] = 4;
        weight_rom[2091] = 5;
        weight_rom[2092] = 5;
        weight_rom[2093] = -7;
        weight_rom[2094] = -10;
        weight_rom[2095] = -16;
        weight_rom[2096] = -53;
        weight_rom[2097] = -69;
        weight_rom[2098] = -23;
        weight_rom[2099] = -6;
        weight_rom[2100] = 3;
        weight_rom[2101] = 12;
        weight_rom[2102] = 7;
        weight_rom[2103] = 21;
        weight_rom[2104] = -10;
        weight_rom[2105] = 8;
        weight_rom[2106] = -14;
        weight_rom[2107] = -26;
        weight_rom[2108] = -19;
        weight_rom[2109] = -28;
        weight_rom[2110] = -28;
        weight_rom[2111] = -35;
        weight_rom[2112] = -31;
        weight_rom[2113] = -31;
        weight_rom[2114] = -20;
        weight_rom[2115] = -12;
        weight_rom[2116] = 0;
        weight_rom[2117] = 12;
        weight_rom[2118] = 9;
        weight_rom[2119] = 7;
        weight_rom[2120] = -8;
        weight_rom[2121] = -2;
        weight_rom[2122] = -15;
        weight_rom[2123] = -2;
        weight_rom[2124] = -38;
        weight_rom[2125] = -55;
        weight_rom[2126] = -24;
        weight_rom[2127] = -4;
        weight_rom[2128] = 2;
        weight_rom[2129] = -11;
        weight_rom[2130] = 5;
        weight_rom[2131] = -8;
        weight_rom[2132] = -3;
        weight_rom[2133] = -2;
        weight_rom[2134] = -8;
        weight_rom[2135] = -15;
        weight_rom[2136] = -30;
        weight_rom[2137] = -22;
        weight_rom[2138] = -29;
        weight_rom[2139] = -35;
        weight_rom[2140] = -38;
        weight_rom[2141] = -25;
        weight_rom[2142] = -15;
        weight_rom[2143] = 1;
        weight_rom[2144] = -2;
        weight_rom[2145] = 6;
        weight_rom[2146] = -2;
        weight_rom[2147] = 3;
        weight_rom[2148] = 8;
        weight_rom[2149] = -9;
        weight_rom[2150] = -8;
        weight_rom[2151] = -27;
        weight_rom[2152] = -33;
        weight_rom[2153] = -18;
        weight_rom[2154] = -20;
        weight_rom[2155] = 1;
        weight_rom[2156] = -4;
        weight_rom[2157] = -3;
        weight_rom[2158] = -6;
        weight_rom[2159] = -31;
        weight_rom[2160] = -13;
        weight_rom[2161] = -17;
        weight_rom[2162] = -12;
        weight_rom[2163] = -12;
        weight_rom[2164] = -18;
        weight_rom[2165] = -23;
        weight_rom[2166] = -26;
        weight_rom[2167] = -27;
        weight_rom[2168] = -26;
        weight_rom[2169] = -16;
        weight_rom[2170] = -11;
        weight_rom[2171] = -6;
        weight_rom[2172] = 1;
        weight_rom[2173] = -1;
        weight_rom[2174] = -11;
        weight_rom[2175] = -3;
        weight_rom[2176] = -8;
        weight_rom[2177] = -11;
        weight_rom[2178] = -7;
        weight_rom[2179] = -36;
        weight_rom[2180] = -31;
        weight_rom[2181] = -27;
        weight_rom[2182] = -19;
        weight_rom[2183] = -3;
        weight_rom[2184] = -4;
        weight_rom[2185] = -3;
        weight_rom[2186] = -6;
        weight_rom[2187] = -7;
        weight_rom[2188] = -11;
        weight_rom[2189] = -26;
        weight_rom[2190] = -29;
        weight_rom[2191] = -5;
        weight_rom[2192] = -13;
        weight_rom[2193] = -19;
        weight_rom[2194] = -16;
        weight_rom[2195] = -7;
        weight_rom[2196] = 0;
        weight_rom[2197] = 4;
        weight_rom[2198] = -3;
        weight_rom[2199] = 2;
        weight_rom[2200] = -1;
        weight_rom[2201] = -7;
        weight_rom[2202] = -14;
        weight_rom[2203] = -5;
        weight_rom[2204] = -15;
        weight_rom[2205] = -8;
        weight_rom[2206] = -4;
        weight_rom[2207] = 4;
        weight_rom[2208] = -20;
        weight_rom[2209] = -17;
        weight_rom[2210] = -9;
        weight_rom[2211] = 3;
        weight_rom[2212] = -2;
        weight_rom[2213] = -4;
        weight_rom[2214] = 19;
        weight_rom[2215] = 32;
        weight_rom[2216] = 10;
        weight_rom[2217] = -21;
        weight_rom[2218] = -10;
        weight_rom[2219] = 3;
        weight_rom[2220] = 1;
        weight_rom[2221] = -3;
        weight_rom[2222] = 3;
        weight_rom[2223] = 0;
        weight_rom[2224] = -4;
        weight_rom[2225] = 10;
        weight_rom[2226] = 14;
        weight_rom[2227] = -1;
        weight_rom[2228] = 9;
        weight_rom[2229] = 4;
        weight_rom[2230] = 4;
        weight_rom[2231] = 2;
        weight_rom[2232] = 2;
        weight_rom[2233] = 12;
        weight_rom[2234] = -1;
        weight_rom[2235] = 7;
        weight_rom[2236] = -9;
        weight_rom[2237] = -25;
        weight_rom[2238] = -10;
        weight_rom[2239] = 1;
        weight_rom[2240] = -1;
        weight_rom[2241] = -4;
        weight_rom[2242] = 9;
        weight_rom[2243] = 35;
        weight_rom[2244] = 32;
        weight_rom[2245] = 13;
        weight_rom[2246] = 9;
        weight_rom[2247] = 33;
        weight_rom[2248] = 32;
        weight_rom[2249] = 10;
        weight_rom[2250] = 28;
        weight_rom[2251] = 29;
        weight_rom[2252] = 12;
        weight_rom[2253] = 11;
        weight_rom[2254] = 14;
        weight_rom[2255] = 14;
        weight_rom[2256] = 34;
        weight_rom[2257] = 3;
        weight_rom[2258] = 21;
        weight_rom[2259] = 33;
        weight_rom[2260] = 23;
        weight_rom[2261] = 19;
        weight_rom[2262] = 13;
        weight_rom[2263] = 16;
        weight_rom[2264] = -13;
        weight_rom[2265] = -28;
        weight_rom[2266] = 4;
        weight_rom[2267] = -2;
        weight_rom[2268] = -1;
        weight_rom[2269] = -2;
        weight_rom[2270] = -1;
        weight_rom[2271] = -13;
        weight_rom[2272] = 15;
        weight_rom[2273] = 46;
        weight_rom[2274] = 38;
        weight_rom[2275] = 59;
        weight_rom[2276] = 49;
        weight_rom[2277] = 56;
        weight_rom[2278] = 73;
        weight_rom[2279] = 62;
        weight_rom[2280] = 44;
        weight_rom[2281] = 47;
        weight_rom[2282] = 46;
        weight_rom[2283] = 44;
        weight_rom[2284] = 42;
        weight_rom[2285] = 32;
        weight_rom[2286] = 36;
        weight_rom[2287] = 46;
        weight_rom[2288] = 40;
        weight_rom[2289] = 28;
        weight_rom[2290] = 8;
        weight_rom[2291] = -4;
        weight_rom[2292] = -8;
        weight_rom[2293] = 3;
        weight_rom[2294] = 3;
        weight_rom[2295] = 0;
        weight_rom[2296] = 4;
        weight_rom[2297] = -2;
        weight_rom[2298] = 1;
        weight_rom[2299] = 3;
        weight_rom[2300] = 27;
        weight_rom[2301] = 26;
        weight_rom[2302] = 36;
        weight_rom[2303] = 47;
        weight_rom[2304] = 37;
        weight_rom[2305] = 31;
        weight_rom[2306] = 27;
        weight_rom[2307] = 21;
        weight_rom[2308] = 15;
        weight_rom[2309] = 37;
        weight_rom[2310] = 39;
        weight_rom[2311] = 6;
        weight_rom[2312] = 27;
        weight_rom[2313] = 31;
        weight_rom[2314] = 38;
        weight_rom[2315] = 12;
        weight_rom[2316] = 16;
        weight_rom[2317] = 23;
        weight_rom[2318] = 8;
        weight_rom[2319] = 10;
        weight_rom[2320] = -4;
        weight_rom[2321] = -2;
        weight_rom[2322] = -3;
        weight_rom[2323] = 2;
        weight_rom[2324] = -3;
        weight_rom[2325] = -1;
        weight_rom[2326] = -1;
        weight_rom[2327] = 3;
        weight_rom[2328] = 2;
        weight_rom[2329] = -23;
        weight_rom[2330] = -38;
        weight_rom[2331] = 8;
        weight_rom[2332] = -5;
        weight_rom[2333] = -5;
        weight_rom[2334] = -6;
        weight_rom[2335] = 1;
        weight_rom[2336] = 1;
        weight_rom[2337] = -39;
        weight_rom[2338] = 4;
        weight_rom[2339] = 2;
        weight_rom[2340] = 0;
        weight_rom[2341] = -28;
        weight_rom[2342] = 5;
        weight_rom[2343] = 13;
        weight_rom[2344] = 4;
        weight_rom[2345] = 3;
        weight_rom[2346] = 19;
        weight_rom[2347] = 3;
        weight_rom[2348] = 4;
        weight_rom[2349] = 1;
        weight_rom[2350] = -1;
        weight_rom[2351] = -4;
        weight_rom[2352] = -3;
        weight_rom[2353] = 1;
        weight_rom[2354] = -1;
        weight_rom[2355] = 0;
        weight_rom[2356] = 1;
        weight_rom[2357] = -2;
        weight_rom[2358] = -4;
        weight_rom[2359] = 0;
        weight_rom[2360] = -1;
        weight_rom[2361] = 1;
        weight_rom[2362] = 4;
        weight_rom[2363] = 0;
        weight_rom[2364] = 1;
        weight_rom[2365] = 14;
        weight_rom[2366] = 4;
        weight_rom[2367] = -4;
        weight_rom[2368] = -4;
        weight_rom[2369] = -5;
        weight_rom[2370] = -2;
        weight_rom[2371] = -4;
        weight_rom[2372] = 2;
        weight_rom[2373] = 0;
        weight_rom[2374] = 1;
        weight_rom[2375] = -2;
        weight_rom[2376] = 3;
        weight_rom[2377] = 1;
        weight_rom[2378] = -3;
        weight_rom[2379] = 3;
        weight_rom[2380] = -2;
        weight_rom[2381] = -2;
        weight_rom[2382] = 1;
        weight_rom[2383] = -4;
        weight_rom[2384] = -1;
        weight_rom[2385] = 1;
        weight_rom[2386] = 3;
        weight_rom[2387] = 4;
        weight_rom[2388] = -13;
        weight_rom[2389] = 7;
        weight_rom[2390] = 17;
        weight_rom[2391] = 6;
        weight_rom[2392] = 16;
        weight_rom[2393] = 38;
        weight_rom[2394] = -1;
        weight_rom[2395] = -2;
        weight_rom[2396] = -40;
        weight_rom[2397] = 3;
        weight_rom[2398] = 36;
        weight_rom[2399] = 22;
        weight_rom[2400] = 26;
        weight_rom[2401] = 19;
        weight_rom[2402] = 14;
        weight_rom[2403] = 13;
        weight_rom[2404] = -4;
        weight_rom[2405] = -1;
        weight_rom[2406] = 2;
        weight_rom[2407] = -3;
        weight_rom[2408] = -2;
        weight_rom[2409] = 3;
        weight_rom[2410] = -3;
        weight_rom[2411] = -2;
        weight_rom[2412] = 16;
        weight_rom[2413] = 2;
        weight_rom[2414] = 0;
        weight_rom[2415] = 4;
        weight_rom[2416] = -2;
        weight_rom[2417] = -1;
        weight_rom[2418] = 11;
        weight_rom[2419] = -13;
        weight_rom[2420] = 1;
        weight_rom[2421] = -4;
        weight_rom[2422] = -14;
        weight_rom[2423] = 0;
        weight_rom[2424] = -6;
        weight_rom[2425] = 3;
        weight_rom[2426] = 14;
        weight_rom[2427] = 19;
        weight_rom[2428] = 26;
        weight_rom[2429] = 13;
        weight_rom[2430] = 39;
        weight_rom[2431] = 23;
        weight_rom[2432] = -5;
        weight_rom[2433] = -13;
        weight_rom[2434] = 0;
        weight_rom[2435] = -3;
        weight_rom[2436] = -2;
        weight_rom[2437] = 1;
        weight_rom[2438] = 4;
        weight_rom[2439] = -1;
        weight_rom[2440] = 2;
        weight_rom[2441] = 4;
        weight_rom[2442] = -9;
        weight_rom[2443] = -7;
        weight_rom[2444] = -10;
        weight_rom[2445] = -33;
        weight_rom[2446] = -7;
        weight_rom[2447] = -13;
        weight_rom[2448] = -21;
        weight_rom[2449] = -26;
        weight_rom[2450] = -29;
        weight_rom[2451] = -15;
        weight_rom[2452] = -18;
        weight_rom[2453] = -14;
        weight_rom[2454] = -6;
        weight_rom[2455] = 16;
        weight_rom[2456] = 12;
        weight_rom[2457] = 19;
        weight_rom[2458] = 10;
        weight_rom[2459] = 12;
        weight_rom[2460] = 3;
        weight_rom[2461] = -24;
        weight_rom[2462] = -2;
        weight_rom[2463] = -1;
        weight_rom[2464] = -2;
        weight_rom[2465] = -4;
        weight_rom[2466] = 11;
        weight_rom[2467] = 1;
        weight_rom[2468] = 8;
        weight_rom[2469] = 0;
        weight_rom[2470] = -37;
        weight_rom[2471] = -24;
        weight_rom[2472] = -44;
        weight_rom[2473] = -51;
        weight_rom[2474] = -36;
        weight_rom[2475] = -28;
        weight_rom[2476] = -40;
        weight_rom[2477] = -17;
        weight_rom[2478] = -28;
        weight_rom[2479] = -24;
        weight_rom[2480] = -19;
        weight_rom[2481] = -12;
        weight_rom[2482] = -12;
        weight_rom[2483] = 6;
        weight_rom[2484] = -3;
        weight_rom[2485] = 9;
        weight_rom[2486] = 16;
        weight_rom[2487] = 34;
        weight_rom[2488] = -5;
        weight_rom[2489] = -21;
        weight_rom[2490] = -20;
        weight_rom[2491] = 4;
        weight_rom[2492] = -2;
        weight_rom[2493] = 1;
        weight_rom[2494] = 1;
        weight_rom[2495] = 1;
        weight_rom[2496] = 23;
        weight_rom[2497] = -9;
        weight_rom[2498] = -29;
        weight_rom[2499] = -39;
        weight_rom[2500] = -56;
        weight_rom[2501] = -36;
        weight_rom[2502] = -22;
        weight_rom[2503] = -44;
        weight_rom[2504] = -22;
        weight_rom[2505] = -17;
        weight_rom[2506] = -15;
        weight_rom[2507] = -2;
        weight_rom[2508] = 4;
        weight_rom[2509] = -7;
        weight_rom[2510] = 2;
        weight_rom[2511] = 16;
        weight_rom[2512] = 3;
        weight_rom[2513] = 15;
        weight_rom[2514] = 9;
        weight_rom[2515] = 24;
        weight_rom[2516] = 21;
        weight_rom[2517] = -17;
        weight_rom[2518] = 4;
        weight_rom[2519] = 2;
        weight_rom[2520] = -4;
        weight_rom[2521] = -3;
        weight_rom[2522] = 0;
        weight_rom[2523] = 14;
        weight_rom[2524] = -1;
        weight_rom[2525] = -23;
        weight_rom[2526] = -38;
        weight_rom[2527] = -50;
        weight_rom[2528] = -50;
        weight_rom[2529] = -33;
        weight_rom[2530] = -22;
        weight_rom[2531] = -15;
        weight_rom[2532] = -8;
        weight_rom[2533] = -9;
        weight_rom[2534] = -5;
        weight_rom[2535] = -6;
        weight_rom[2536] = -6;
        weight_rom[2537] = -5;
        weight_rom[2538] = -2;
        weight_rom[2539] = 3;
        weight_rom[2540] = 9;
        weight_rom[2541] = 8;
        weight_rom[2542] = 13;
        weight_rom[2543] = 29;
        weight_rom[2544] = 32;
        weight_rom[2545] = -1;
        weight_rom[2546] = 12;
        weight_rom[2547] = 8;
        weight_rom[2548] = 1;
        weight_rom[2549] = 15;
        weight_rom[2550] = -12;
        weight_rom[2551] = 10;
        weight_rom[2552] = 6;
        weight_rom[2553] = -22;
        weight_rom[2554] = -52;
        weight_rom[2555] = -42;
        weight_rom[2556] = -35;
        weight_rom[2557] = -23;
        weight_rom[2558] = -4;
        weight_rom[2559] = -10;
        weight_rom[2560] = 2;
        weight_rom[2561] = 0;
        weight_rom[2562] = 7;
        weight_rom[2563] = -2;
        weight_rom[2564] = -10;
        weight_rom[2565] = 1;
        weight_rom[2566] = -5;
        weight_rom[2567] = 4;
        weight_rom[2568] = 13;
        weight_rom[2569] = 13;
        weight_rom[2570] = 3;
        weight_rom[2571] = 13;
        weight_rom[2572] = -3;
        weight_rom[2573] = -8;
        weight_rom[2574] = 15;
        weight_rom[2575] = -5;
        weight_rom[2576] = 2;
        weight_rom[2577] = 10;
        weight_rom[2578] = -17;
        weight_rom[2579] = 22;
        weight_rom[2580] = -13;
        weight_rom[2581] = -23;
        weight_rom[2582] = -38;
        weight_rom[2583] = -32;
        weight_rom[2584] = -34;
        weight_rom[2585] = -26;
        weight_rom[2586] = -24;
        weight_rom[2587] = -8;
        weight_rom[2588] = -1;
        weight_rom[2589] = 5;
        weight_rom[2590] = 10;
        weight_rom[2591] = 9;
        weight_rom[2592] = -5;
        weight_rom[2593] = 9;
        weight_rom[2594] = -4;
        weight_rom[2595] = -10;
        weight_rom[2596] = -9;
        weight_rom[2597] = 5;
        weight_rom[2598] = -6;
        weight_rom[2599] = -13;
        weight_rom[2600] = -16;
        weight_rom[2601] = -8;
        weight_rom[2602] = -15;
        weight_rom[2603] = 11;
        weight_rom[2604] = -15;
        weight_rom[2605] = 12;
        weight_rom[2606] = -3;
        weight_rom[2607] = -13;
        weight_rom[2608] = -23;
        weight_rom[2609] = -35;
        weight_rom[2610] = -25;
        weight_rom[2611] = -18;
        weight_rom[2612] = -31;
        weight_rom[2613] = -48;
        weight_rom[2614] = -24;
        weight_rom[2615] = -11;
        weight_rom[2616] = -13;
        weight_rom[2617] = 8;
        weight_rom[2618] = 25;
        weight_rom[2619] = 31;
        weight_rom[2620] = 4;
        weight_rom[2621] = 2;
        weight_rom[2622] = -7;
        weight_rom[2623] = -16;
        weight_rom[2624] = -12;
        weight_rom[2625] = -8;
        weight_rom[2626] = -17;
        weight_rom[2627] = -9;
        weight_rom[2628] = 5;
        weight_rom[2629] = -14;
        weight_rom[2630] = 1;
        weight_rom[2631] = 1;
        weight_rom[2632] = -15;
        weight_rom[2633] = 3;
        weight_rom[2634] = -25;
        weight_rom[2635] = -26;
        weight_rom[2636] = -39;
        weight_rom[2637] = -44;
        weight_rom[2638] = -49;
        weight_rom[2639] = -34;
        weight_rom[2640] = -27;
        weight_rom[2641] = -45;
        weight_rom[2642] = -43;
        weight_rom[2643] = -21;
        weight_rom[2644] = -14;
        weight_rom[2645] = 36;
        weight_rom[2646] = 34;
        weight_rom[2647] = 40;
        weight_rom[2648] = 28;
        weight_rom[2649] = 12;
        weight_rom[2650] = 9;
        weight_rom[2651] = -8;
        weight_rom[2652] = -9;
        weight_rom[2653] = -27;
        weight_rom[2654] = -23;
        weight_rom[2655] = -11;
        weight_rom[2656] = -12;
        weight_rom[2657] = 15;
        weight_rom[2658] = -7;
        weight_rom[2659] = -10;
        weight_rom[2660] = -2;
        weight_rom[2661] = -14;
        weight_rom[2662] = -27;
        weight_rom[2663] = -30;
        weight_rom[2664] = -43;
        weight_rom[2665] = -30;
        weight_rom[2666] = -30;
        weight_rom[2667] = -32;
        weight_rom[2668] = -30;
        weight_rom[2669] = -32;
        weight_rom[2670] = -26;
        weight_rom[2671] = -11;
        weight_rom[2672] = 16;
        weight_rom[2673] = 46;
        weight_rom[2674] = 51;
        weight_rom[2675] = 30;
        weight_rom[2676] = 22;
        weight_rom[2677] = -4;
        weight_rom[2678] = -11;
        weight_rom[2679] = -14;
        weight_rom[2680] = -15;
        weight_rom[2681] = -16;
        weight_rom[2682] = -43;
        weight_rom[2683] = -20;
        weight_rom[2684] = -24;
        weight_rom[2685] = -29;
        weight_rom[2686] = -20;
        weight_rom[2687] = 4;
        weight_rom[2688] = -2;
        weight_rom[2689] = -14;
        weight_rom[2690] = -24;
        weight_rom[2691] = -34;
        weight_rom[2692] = -36;
        weight_rom[2693] = -43;
        weight_rom[2694] = -14;
        weight_rom[2695] = -22;
        weight_rom[2696] = -19;
        weight_rom[2697] = -14;
        weight_rom[2698] = 3;
        weight_rom[2699] = 13;
        weight_rom[2700] = 33;
        weight_rom[2701] = 50;
        weight_rom[2702] = 42;
        weight_rom[2703] = 27;
        weight_rom[2704] = 4;
        weight_rom[2705] = -2;
        weight_rom[2706] = -3;
        weight_rom[2707] = -23;
        weight_rom[2708] = -18;
        weight_rom[2709] = -23;
        weight_rom[2710] = -50;
        weight_rom[2711] = -39;
        weight_rom[2712] = -50;
        weight_rom[2713] = -45;
        weight_rom[2714] = -43;
        weight_rom[2715] = 3;
        weight_rom[2716] = 2;
        weight_rom[2717] = -4;
        weight_rom[2718] = -11;
        weight_rom[2719] = -20;
        weight_rom[2720] = -22;
        weight_rom[2721] = -22;
        weight_rom[2722] = -11;
        weight_rom[2723] = -20;
        weight_rom[2724] = -14;
        weight_rom[2725] = 4;
        weight_rom[2726] = 18;
        weight_rom[2727] = 15;
        weight_rom[2728] = 34;
        weight_rom[2729] = 33;
        weight_rom[2730] = 25;
        weight_rom[2731] = 23;
        weight_rom[2732] = -6;
        weight_rom[2733] = 7;
        weight_rom[2734] = 5;
        weight_rom[2735] = -5;
        weight_rom[2736] = 8;
        weight_rom[2737] = -3;
        weight_rom[2738] = -41;
        weight_rom[2739] = -65;
        weight_rom[2740] = -73;
        weight_rom[2741] = -60;
        weight_rom[2742] = -26;
        weight_rom[2743] = -15;
        weight_rom[2744] = 4;
        weight_rom[2745] = -4;
        weight_rom[2746] = -15;
        weight_rom[2747] = 17;
        weight_rom[2748] = -12;
        weight_rom[2749] = -21;
        weight_rom[2750] = -21;
        weight_rom[2751] = -40;
        weight_rom[2752] = -8;
        weight_rom[2753] = 17;
        weight_rom[2754] = 19;
        weight_rom[2755] = 23;
        weight_rom[2756] = 31;
        weight_rom[2757] = 18;
        weight_rom[2758] = 22;
        weight_rom[2759] = 10;
        weight_rom[2760] = 5;
        weight_rom[2761] = -9;
        weight_rom[2762] = 0;
        weight_rom[2763] = 2;
        weight_rom[2764] = 13;
        weight_rom[2765] = -10;
        weight_rom[2766] = -33;
        weight_rom[2767] = -76;
        weight_rom[2768] = -77;
        weight_rom[2769] = -60;
        weight_rom[2770] = -30;
        weight_rom[2771] = 3;
        weight_rom[2772] = -4;
        weight_rom[2773] = 1;
        weight_rom[2774] = -11;
        weight_rom[2775] = -9;
        weight_rom[2776] = -27;
        weight_rom[2777] = -28;
        weight_rom[2778] = -33;
        weight_rom[2779] = -26;
        weight_rom[2780] = 3;
        weight_rom[2781] = 6;
        weight_rom[2782] = 5;
        weight_rom[2783] = 21;
        weight_rom[2784] = 29;
        weight_rom[2785] = 15;
        weight_rom[2786] = 26;
        weight_rom[2787] = -1;
        weight_rom[2788] = -8;
        weight_rom[2789] = 5;
        weight_rom[2790] = 20;
        weight_rom[2791] = 21;
        weight_rom[2792] = 20;
        weight_rom[2793] = 0;
        weight_rom[2794] = -37;
        weight_rom[2795] = -60;
        weight_rom[2796] = -73;
        weight_rom[2797] = -61;
        weight_rom[2798] = -34;
        weight_rom[2799] = -21;
        weight_rom[2800] = 1;
        weight_rom[2801] = 4;
        weight_rom[2802] = 19;
        weight_rom[2803] = -24;
        weight_rom[2804] = -1;
        weight_rom[2805] = -9;
        weight_rom[2806] = -33;
        weight_rom[2807] = -31;
        weight_rom[2808] = -10;
        weight_rom[2809] = -5;
        weight_rom[2810] = 4;
        weight_rom[2811] = 18;
        weight_rom[2812] = 3;
        weight_rom[2813] = 15;
        weight_rom[2814] = 23;
        weight_rom[2815] = -1;
        weight_rom[2816] = -3;
        weight_rom[2817] = -7;
        weight_rom[2818] = 17;
        weight_rom[2819] = 28;
        weight_rom[2820] = 17;
        weight_rom[2821] = -10;
        weight_rom[2822] = -55;
        weight_rom[2823] = -68;
        weight_rom[2824] = -51;
        weight_rom[2825] = -55;
        weight_rom[2826] = -22;
        weight_rom[2827] = -6;
        weight_rom[2828] = 3;
        weight_rom[2829] = 5;
        weight_rom[2830] = -19;
        weight_rom[2831] = -20;
        weight_rom[2832] = 13;
        weight_rom[2833] = -4;
        weight_rom[2834] = -17;
        weight_rom[2835] = -25;
        weight_rom[2836] = -23;
        weight_rom[2837] = -5;
        weight_rom[2838] = 7;
        weight_rom[2839] = 5;
        weight_rom[2840] = 3;
        weight_rom[2841] = 18;
        weight_rom[2842] = 13;
        weight_rom[2843] = -10;
        weight_rom[2844] = -10;
        weight_rom[2845] = -3;
        weight_rom[2846] = 16;
        weight_rom[2847] = 11;
        weight_rom[2848] = 2;
        weight_rom[2849] = -17;
        weight_rom[2850] = -49;
        weight_rom[2851] = -62;
        weight_rom[2852] = -68;
        weight_rom[2853] = -44;
        weight_rom[2854] = -22;
        weight_rom[2855] = 1;
        weight_rom[2856] = -3;
        weight_rom[2857] = -1;
        weight_rom[2858] = 3;
        weight_rom[2859] = 7;
        weight_rom[2860] = 11;
        weight_rom[2861] = -1;
        weight_rom[2862] = -11;
        weight_rom[2863] = -21;
        weight_rom[2864] = -20;
        weight_rom[2865] = -16;
        weight_rom[2866] = -15;
        weight_rom[2867] = 3;
        weight_rom[2868] = 25;
        weight_rom[2869] = 14;
        weight_rom[2870] = 20;
        weight_rom[2871] = 2;
        weight_rom[2872] = -1;
        weight_rom[2873] = 4;
        weight_rom[2874] = 21;
        weight_rom[2875] = -8;
        weight_rom[2876] = -12;
        weight_rom[2877] = -24;
        weight_rom[2878] = -59;
        weight_rom[2879] = -59;
        weight_rom[2880] = -57;
        weight_rom[2881] = -32;
        weight_rom[2882] = 2;
        weight_rom[2883] = -3;
        weight_rom[2884] = 0;
        weight_rom[2885] = -3;
        weight_rom[2886] = 6;
        weight_rom[2887] = 13;
        weight_rom[2888] = 1;
        weight_rom[2889] = -11;
        weight_rom[2890] = 6;
        weight_rom[2891] = -6;
        weight_rom[2892] = -21;
        weight_rom[2893] = -2;
        weight_rom[2894] = -5;
        weight_rom[2895] = 23;
        weight_rom[2896] = 26;
        weight_rom[2897] = 17;
        weight_rom[2898] = 13;
        weight_rom[2899] = 21;
        weight_rom[2900] = 27;
        weight_rom[2901] = 6;
        weight_rom[2902] = 14;
        weight_rom[2903] = -2;
        weight_rom[2904] = -18;
        weight_rom[2905] = -42;
        weight_rom[2906] = -76;
        weight_rom[2907] = -67;
        weight_rom[2908] = -27;
        weight_rom[2909] = -15;
        weight_rom[2910] = 0;
        weight_rom[2911] = -3;
        weight_rom[2912] = 3;
        weight_rom[2913] = -5;
        weight_rom[2914] = -1;
        weight_rom[2915] = 4;
        weight_rom[2916] = -2;
        weight_rom[2917] = -9;
        weight_rom[2918] = 3;
        weight_rom[2919] = 0;
        weight_rom[2920] = 1;
        weight_rom[2921] = 0;
        weight_rom[2922] = 4;
        weight_rom[2923] = 7;
        weight_rom[2924] = 6;
        weight_rom[2925] = 10;
        weight_rom[2926] = 26;
        weight_rom[2927] = 17;
        weight_rom[2928] = 17;
        weight_rom[2929] = 13;
        weight_rom[2930] = 6;
        weight_rom[2931] = -15;
        weight_rom[2932] = -31;
        weight_rom[2933] = -34;
        weight_rom[2934] = -68;
        weight_rom[2935] = -39;
        weight_rom[2936] = -21;
        weight_rom[2937] = -1;
        weight_rom[2938] = 10;
        weight_rom[2939] = 4;
        weight_rom[2940] = 5;
        weight_rom[2941] = -4;
        weight_rom[2942] = 2;
        weight_rom[2943] = 2;
        weight_rom[2944] = -6;
        weight_rom[2945] = 4;
        weight_rom[2946] = -2;
        weight_rom[2947] = 8;
        weight_rom[2948] = 11;
        weight_rom[2949] = 3;
        weight_rom[2950] = 11;
        weight_rom[2951] = 1;
        weight_rom[2952] = 7;
        weight_rom[2953] = 19;
        weight_rom[2954] = 25;
        weight_rom[2955] = 23;
        weight_rom[2956] = 13;
        weight_rom[2957] = -2;
        weight_rom[2958] = -12;
        weight_rom[2959] = -32;
        weight_rom[2960] = -32;
        weight_rom[2961] = -42;
        weight_rom[2962] = -65;
        weight_rom[2963] = -34;
        weight_rom[2964] = -4;
        weight_rom[2965] = -7;
        weight_rom[2966] = 15;
        weight_rom[2967] = 1;
        weight_rom[2968] = -4;
        weight_rom[2969] = 0;
        weight_rom[2970] = 16;
        weight_rom[2971] = -3;
        weight_rom[2972] = 0;
        weight_rom[2973] = 32;
        weight_rom[2974] = 17;
        weight_rom[2975] = 4;
        weight_rom[2976] = 5;
        weight_rom[2977] = 7;
        weight_rom[2978] = 11;
        weight_rom[2979] = 7;
        weight_rom[2980] = 12;
        weight_rom[2981] = 7;
        weight_rom[2982] = 28;
        weight_rom[2983] = 18;
        weight_rom[2984] = 10;
        weight_rom[2985] = 6;
        weight_rom[2986] = -21;
        weight_rom[2987] = -27;
        weight_rom[2988] = -45;
        weight_rom[2989] = -34;
        weight_rom[2990] = -29;
        weight_rom[2991] = -14;
        weight_rom[2992] = -8;
        weight_rom[2993] = 1;
        weight_rom[2994] = 9;
        weight_rom[2995] = -3;
        weight_rom[2996] = -2;
        weight_rom[2997] = 2;
        weight_rom[2998] = 1;
        weight_rom[2999] = -13;
        weight_rom[3000] = 7;
        weight_rom[3001] = 27;
        weight_rom[3002] = 29;
        weight_rom[3003] = 11;
        weight_rom[3004] = 6;
        weight_rom[3005] = 15;
        weight_rom[3006] = 1;
        weight_rom[3007] = 15;
        weight_rom[3008] = 6;
        weight_rom[3009] = 0;
        weight_rom[3010] = -2;
        weight_rom[3011] = 17;
        weight_rom[3012] = -5;
        weight_rom[3013] = -13;
        weight_rom[3014] = -25;
        weight_rom[3015] = -21;
        weight_rom[3016] = -34;
        weight_rom[3017] = -35;
        weight_rom[3018] = -20;
        weight_rom[3019] = -29;
        weight_rom[3020] = 2;
        weight_rom[3021] = 4;
        weight_rom[3022] = 8;
        weight_rom[3023] = 0;
        weight_rom[3024] = 3;
        weight_rom[3025] = 2;
        weight_rom[3026] = 2;
        weight_rom[3027] = -10;
        weight_rom[3028] = -5;
        weight_rom[3029] = -6;
        weight_rom[3030] = 4;
        weight_rom[3031] = -10;
        weight_rom[3032] = -9;
        weight_rom[3033] = 8;
        weight_rom[3034] = -2;
        weight_rom[3035] = -5;
        weight_rom[3036] = -9;
        weight_rom[3037] = -23;
        weight_rom[3038] = -11;
        weight_rom[3039] = -23;
        weight_rom[3040] = -35;
        weight_rom[3041] = -17;
        weight_rom[3042] = -18;
        weight_rom[3043] = 9;
        weight_rom[3044] = -15;
        weight_rom[3045] = -17;
        weight_rom[3046] = 3;
        weight_rom[3047] = -7;
        weight_rom[3048] = -4;
        weight_rom[3049] = 1;
        weight_rom[3050] = -3;
        weight_rom[3051] = -1;
        weight_rom[3052] = 4;
        weight_rom[3053] = 4;
        weight_rom[3054] = -3;
        weight_rom[3055] = 3;
        weight_rom[3056] = -17;
        weight_rom[3057] = -38;
        weight_rom[3058] = -27;
        weight_rom[3059] = -41;
        weight_rom[3060] = -39;
        weight_rom[3061] = -34;
        weight_rom[3062] = -41;
        weight_rom[3063] = -42;
        weight_rom[3064] = -51;
        weight_rom[3065] = -56;
        weight_rom[3066] = -57;
        weight_rom[3067] = -74;
        weight_rom[3068] = -58;
        weight_rom[3069] = -59;
        weight_rom[3070] = -39;
        weight_rom[3071] = -32;
        weight_rom[3072] = 0;
        weight_rom[3073] = -17;
        weight_rom[3074] = -5;
        weight_rom[3075] = 10;
        weight_rom[3076] = -1;
        weight_rom[3077] = 3;
        weight_rom[3078] = 2;
        weight_rom[3079] = 4;
        weight_rom[3080] = 2;
        weight_rom[3081] = 1;
        weight_rom[3082] = 1;
        weight_rom[3083] = 2;
        weight_rom[3084] = -18;
        weight_rom[3085] = -17;
        weight_rom[3086] = -30;
        weight_rom[3087] = -38;
        weight_rom[3088] = -49;
        weight_rom[3089] = -54;
        weight_rom[3090] = -52;
        weight_rom[3091] = -45;
        weight_rom[3092] = -72;
        weight_rom[3093] = -86;
        weight_rom[3094] = -79;
        weight_rom[3095] = -44;
        weight_rom[3096] = -67;
        weight_rom[3097] = -66;
        weight_rom[3098] = -53;
        weight_rom[3099] = -42;
        weight_rom[3100] = -18;
        weight_rom[3101] = -8;
        weight_rom[3102] = -17;
        weight_rom[3103] = -4;
        weight_rom[3104] = -2;
        weight_rom[3105] = 4;
        weight_rom[3106] = 3;
        weight_rom[3107] = -1;
        weight_rom[3108] = 2;
        weight_rom[3109] = -4;
        weight_rom[3110] = 3;
        weight_rom[3111] = -1;
        weight_rom[3112] = -3;
        weight_rom[3113] = 2;
        weight_rom[3114] = 6;
        weight_rom[3115] = -13;
        weight_rom[3116] = -14;
        weight_rom[3117] = -19;
        weight_rom[3118] = -28;
        weight_rom[3119] = -15;
        weight_rom[3120] = -23;
        weight_rom[3121] = -9;
        weight_rom[3122] = -32;
        weight_rom[3123] = -21;
        weight_rom[3124] = -16;
        weight_rom[3125] = -1;
        weight_rom[3126] = -18;
        weight_rom[3127] = -10;
        weight_rom[3128] = 1;
        weight_rom[3129] = 0;
        weight_rom[3130] = -1;
        weight_rom[3131] = 4;
        weight_rom[3132] = 4;
        weight_rom[3133] = 4;
        weight_rom[3134] = -1;
        weight_rom[3135] = 4;
        weight_rom[3136] = 0;
        weight_rom[3137] = 0;
        weight_rom[3138] = -2;
        weight_rom[3139] = -4;
        weight_rom[3140] = -3;
        weight_rom[3141] = 1;
        weight_rom[3142] = 4;
        weight_rom[3143] = -1;
        weight_rom[3144] = -2;
        weight_rom[3145] = 4;
        weight_rom[3146] = -4;
        weight_rom[3147] = 3;
        weight_rom[3148] = 1;
        weight_rom[3149] = -2;
        weight_rom[3150] = 2;
        weight_rom[3151] = -3;
        weight_rom[3152] = -3;
        weight_rom[3153] = -1;
        weight_rom[3154] = 4;
        weight_rom[3155] = 1;
        weight_rom[3156] = 0;
        weight_rom[3157] = -3;
        weight_rom[3158] = 2;
        weight_rom[3159] = 4;
        weight_rom[3160] = 1;
        weight_rom[3161] = -3;
        weight_rom[3162] = -1;
        weight_rom[3163] = 0;
        weight_rom[3164] = -1;
        weight_rom[3165] = -2;
        weight_rom[3166] = 4;
        weight_rom[3167] = -2;
        weight_rom[3168] = -2;
        weight_rom[3169] = 0;
        weight_rom[3170] = 4;
        weight_rom[3171] = -6;
        weight_rom[3172] = -7;
        weight_rom[3173] = -12;
        weight_rom[3174] = -9;
        weight_rom[3175] = -12;
        weight_rom[3176] = -22;
        weight_rom[3177] = -5;
        weight_rom[3178] = -18;
        weight_rom[3179] = -10;
        weight_rom[3180] = -30;
        weight_rom[3181] = -7;
        weight_rom[3182] = -1;
        weight_rom[3183] = -14;
        weight_rom[3184] = -11;
        weight_rom[3185] = -17;
        weight_rom[3186] = -14;
        weight_rom[3187] = -6;
        weight_rom[3188] = 4;
        weight_rom[3189] = 0;
        weight_rom[3190] = -3;
        weight_rom[3191] = -1;
        weight_rom[3192] = -4;
        weight_rom[3193] = 1;
        weight_rom[3194] = 0;
        weight_rom[3195] = -1;
        weight_rom[3196] = -3;
        weight_rom[3197] = 1;
        weight_rom[3198] = -10;
        weight_rom[3199] = -11;
        weight_rom[3200] = -11;
        weight_rom[3201] = -24;
        weight_rom[3202] = -37;
        weight_rom[3203] = -19;
        weight_rom[3204] = -39;
        weight_rom[3205] = -27;
        weight_rom[3206] = -41;
        weight_rom[3207] = -36;
        weight_rom[3208] = -45;
        weight_rom[3209] = -36;
        weight_rom[3210] = -18;
        weight_rom[3211] = -28;
        weight_rom[3212] = -15;
        weight_rom[3213] = -21;
        weight_rom[3214] = -18;
        weight_rom[3215] = -5;
        weight_rom[3216] = -17;
        weight_rom[3217] = -11;
        weight_rom[3218] = 0;
        weight_rom[3219] = 1;
        weight_rom[3220] = 2;
        weight_rom[3221] = 2;
        weight_rom[3222] = 0;
        weight_rom[3223] = -4;
        weight_rom[3224] = -4;
        weight_rom[3225] = 10;
        weight_rom[3226] = -16;
        weight_rom[3227] = -14;
        weight_rom[3228] = -35;
        weight_rom[3229] = -34;
        weight_rom[3230] = -44;
        weight_rom[3231] = -55;
        weight_rom[3232] = -52;
        weight_rom[3233] = -47;
        weight_rom[3234] = -42;
        weight_rom[3235] = -40;
        weight_rom[3236] = -24;
        weight_rom[3237] = -30;
        weight_rom[3238] = -20;
        weight_rom[3239] = -41;
        weight_rom[3240] = -44;
        weight_rom[3241] = -19;
        weight_rom[3242] = -10;
        weight_rom[3243] = -9;
        weight_rom[3244] = -17;
        weight_rom[3245] = -25;
        weight_rom[3246] = 4;
        weight_rom[3247] = -3;
        weight_rom[3248] = 1;
        weight_rom[3249] = 2;
        weight_rom[3250] = 7;
        weight_rom[3251] = -3;
        weight_rom[3252] = 11;
        weight_rom[3253] = -4;
        weight_rom[3254] = 3;
        weight_rom[3255] = -7;
        weight_rom[3256] = -9;
        weight_rom[3257] = 2;
        weight_rom[3258] = 4;
        weight_rom[3259] = -7;
        weight_rom[3260] = 12;
        weight_rom[3261] = 15;
        weight_rom[3262] = 9;
        weight_rom[3263] = 13;
        weight_rom[3264] = 15;
        weight_rom[3265] = 3;
        weight_rom[3266] = 8;
        weight_rom[3267] = 18;
        weight_rom[3268] = 14;
        weight_rom[3269] = -4;
        weight_rom[3270] = -8;
        weight_rom[3271] = -18;
        weight_rom[3272] = -24;
        weight_rom[3273] = -16;
        weight_rom[3274] = 9;
        weight_rom[3275] = -1;
        weight_rom[3276] = -4;
        weight_rom[3277] = -3;
        weight_rom[3278] = 4;
        weight_rom[3279] = 16;
        weight_rom[3280] = 5;
        weight_rom[3281] = 24;
        weight_rom[3282] = 5;
        weight_rom[3283] = 11;
        weight_rom[3284] = 12;
        weight_rom[3285] = -4;
        weight_rom[3286] = -9;
        weight_rom[3287] = 3;
        weight_rom[3288] = 10;
        weight_rom[3289] = 11;
        weight_rom[3290] = 2;
        weight_rom[3291] = 8;
        weight_rom[3292] = 4;
        weight_rom[3293] = 5;
        weight_rom[3294] = 1;
        weight_rom[3295] = 15;
        weight_rom[3296] = 1;
        weight_rom[3297] = 9;
        weight_rom[3298] = -10;
        weight_rom[3299] = -10;
        weight_rom[3300] = 1;
        weight_rom[3301] = -6;
        weight_rom[3302] = -4;
        weight_rom[3303] = -1;
        weight_rom[3304] = -2;
        weight_rom[3305] = -1;
        weight_rom[3306] = -5;
        weight_rom[3307] = -9;
        weight_rom[3308] = -9;
        weight_rom[3309] = -1;
        weight_rom[3310] = -1;
        weight_rom[3311] = 6;
        weight_rom[3312] = -2;
        weight_rom[3313] = -16;
        weight_rom[3314] = -7;
        weight_rom[3315] = -3;
        weight_rom[3316] = -8;
        weight_rom[3317] = -2;
        weight_rom[3318] = -3;
        weight_rom[3319] = 3;
        weight_rom[3320] = 4;
        weight_rom[3321] = 17;
        weight_rom[3322] = 5;
        weight_rom[3323] = 11;
        weight_rom[3324] = 14;
        weight_rom[3325] = 4;
        weight_rom[3326] = -2;
        weight_rom[3327] = -1;
        weight_rom[3328] = -21;
        weight_rom[3329] = 8;
        weight_rom[3330] = -13;
        weight_rom[3331] = -7;
        weight_rom[3332] = 0;
        weight_rom[3333] = -19;
        weight_rom[3334] = -6;
        weight_rom[3335] = 10;
        weight_rom[3336] = 1;
        weight_rom[3337] = -19;
        weight_rom[3338] = -10;
        weight_rom[3339] = -16;
        weight_rom[3340] = -10;
        weight_rom[3341] = -11;
        weight_rom[3342] = -14;
        weight_rom[3343] = -21;
        weight_rom[3344] = -16;
        weight_rom[3345] = -11;
        weight_rom[3346] = -11;
        weight_rom[3347] = -1;
        weight_rom[3348] = 5;
        weight_rom[3349] = 1;
        weight_rom[3350] = 12;
        weight_rom[3351] = 17;
        weight_rom[3352] = 17;
        weight_rom[3353] = 9;
        weight_rom[3354] = -11;
        weight_rom[3355] = -11;
        weight_rom[3356] = -24;
        weight_rom[3357] = -20;
        weight_rom[3358] = -11;
        weight_rom[3359] = 3;
        weight_rom[3360] = 5;
        weight_rom[3361] = -20;
        weight_rom[3362] = -1;
        weight_rom[3363] = -13;
        weight_rom[3364] = -6;
        weight_rom[3365] = -7;
        weight_rom[3366] = 1;
        weight_rom[3367] = -7;
        weight_rom[3368] = -6;
        weight_rom[3369] = -7;
        weight_rom[3370] = -13;
        weight_rom[3371] = -20;
        weight_rom[3372] = -2;
        weight_rom[3373] = 2;
        weight_rom[3374] = -2;
        weight_rom[3375] = -5;
        weight_rom[3376] = -7;
        weight_rom[3377] = -6;
        weight_rom[3378] = 17;
        weight_rom[3379] = 5;
        weight_rom[3380] = -2;
        weight_rom[3381] = 7;
        weight_rom[3382] = -10;
        weight_rom[3383] = -23;
        weight_rom[3384] = -26;
        weight_rom[3385] = -12;
        weight_rom[3386] = 2;
        weight_rom[3387] = 1;
        weight_rom[3388] = -11;
        weight_rom[3389] = -17;
        weight_rom[3390] = -23;
        weight_rom[3391] = -21;
        weight_rom[3392] = -14;
        weight_rom[3393] = -6;
        weight_rom[3394] = 5;
        weight_rom[3395] = -5;
        weight_rom[3396] = -4;
        weight_rom[3397] = -7;
        weight_rom[3398] = -2;
        weight_rom[3399] = 0;
        weight_rom[3400] = 4;
        weight_rom[3401] = 13;
        weight_rom[3402] = 0;
        weight_rom[3403] = 7;
        weight_rom[3404] = 11;
        weight_rom[3405] = 14;
        weight_rom[3406] = 15;
        weight_rom[3407] = 9;
        weight_rom[3408] = 2;
        weight_rom[3409] = -2;
        weight_rom[3410] = -13;
        weight_rom[3411] = -29;
        weight_rom[3412] = -42;
        weight_rom[3413] = -27;
        weight_rom[3414] = 3;
        weight_rom[3415] = -16;
        weight_rom[3416] = -8;
        weight_rom[3417] = -11;
        weight_rom[3418] = -19;
        weight_rom[3419] = -35;
        weight_rom[3420] = -7;
        weight_rom[3421] = -18;
        weight_rom[3422] = -6;
        weight_rom[3423] = -3;
        weight_rom[3424] = 8;
        weight_rom[3425] = 3;
        weight_rom[3426] = 12;
        weight_rom[3427] = 12;
        weight_rom[3428] = 20;
        weight_rom[3429] = 11;
        weight_rom[3430] = 15;
        weight_rom[3431] = 6;
        weight_rom[3432] = 9;
        weight_rom[3433] = 8;
        weight_rom[3434] = 13;
        weight_rom[3435] = 14;
        weight_rom[3436] = 6;
        weight_rom[3437] = -6;
        weight_rom[3438] = -11;
        weight_rom[3439] = -44;
        weight_rom[3440] = -65;
        weight_rom[3441] = -62;
        weight_rom[3442] = -28;
        weight_rom[3443] = 15;
        weight_rom[3444] = 11;
        weight_rom[3445] = -10;
        weight_rom[3446] = -38;
        weight_rom[3447] = -20;
        weight_rom[3448] = -25;
        weight_rom[3449] = -21;
        weight_rom[3450] = -6;
        weight_rom[3451] = 9;
        weight_rom[3452] = 14;
        weight_rom[3453] = 18;
        weight_rom[3454] = 29;
        weight_rom[3455] = 34;
        weight_rom[3456] = 32;
        weight_rom[3457] = 27;
        weight_rom[3458] = 41;
        weight_rom[3459] = 35;
        weight_rom[3460] = 22;
        weight_rom[3461] = 25;
        weight_rom[3462] = 20;
        weight_rom[3463] = 8;
        weight_rom[3464] = 8;
        weight_rom[3465] = 4;
        weight_rom[3466] = -4;
        weight_rom[3467] = -32;
        weight_rom[3468] = -36;
        weight_rom[3469] = -39;
        weight_rom[3470] = -3;
        weight_rom[3471] = 2;
        weight_rom[3472] = 9;
        weight_rom[3473] = -4;
        weight_rom[3474] = -19;
        weight_rom[3475] = -20;
        weight_rom[3476] = -8;
        weight_rom[3477] = -10;
        weight_rom[3478] = -3;
        weight_rom[3479] = 15;
        weight_rom[3480] = 14;
        weight_rom[3481] = 20;
        weight_rom[3482] = 11;
        weight_rom[3483] = 26;
        weight_rom[3484] = 14;
        weight_rom[3485] = 34;
        weight_rom[3486] = 44;
        weight_rom[3487] = 33;
        weight_rom[3488] = 30;
        weight_rom[3489] = 37;
        weight_rom[3490] = 27;
        weight_rom[3491] = 21;
        weight_rom[3492] = 31;
        weight_rom[3493] = 27;
        weight_rom[3494] = 20;
        weight_rom[3495] = 10;
        weight_rom[3496] = -11;
        weight_rom[3497] = -25;
        weight_rom[3498] = -17;
        weight_rom[3499] = -4;
        weight_rom[3500] = -1;
        weight_rom[3501] = -11;
        weight_rom[3502] = -33;
        weight_rom[3503] = -10;
        weight_rom[3504] = -6;
        weight_rom[3505] = -13;
        weight_rom[3506] = -5;
        weight_rom[3507] = 16;
        weight_rom[3508] = 4;
        weight_rom[3509] = 13;
        weight_rom[3510] = 7;
        weight_rom[3511] = -3;
        weight_rom[3512] = 6;
        weight_rom[3513] = 25;
        weight_rom[3514] = 28;
        weight_rom[3515] = 44;
        weight_rom[3516] = 41;
        weight_rom[3517] = 32;
        weight_rom[3518] = 25;
        weight_rom[3519] = 19;
        weight_rom[3520] = 16;
        weight_rom[3521] = 15;
        weight_rom[3522] = -2;
        weight_rom[3523] = -14;
        weight_rom[3524] = -28;
        weight_rom[3525] = -22;
        weight_rom[3526] = -21;
        weight_rom[3527] = -14;
        weight_rom[3528] = 1;
        weight_rom[3529] = -9;
        weight_rom[3530] = -19;
        weight_rom[3531] = -9;
        weight_rom[3532] = -13;
        weight_rom[3533] = -29;
        weight_rom[3534] = -13;
        weight_rom[3535] = -15;
        weight_rom[3536] = -19;
        weight_rom[3537] = -10;
        weight_rom[3538] = -9;
        weight_rom[3539] = -4;
        weight_rom[3540] = 14;
        weight_rom[3541] = 25;
        weight_rom[3542] = 28;
        weight_rom[3543] = 26;
        weight_rom[3544] = 28;
        weight_rom[3545] = 23;
        weight_rom[3546] = 16;
        weight_rom[3547] = -6;
        weight_rom[3548] = -31;
        weight_rom[3549] = -25;
        weight_rom[3550] = -31;
        weight_rom[3551] = -31;
        weight_rom[3552] = -44;
        weight_rom[3553] = -22;
        weight_rom[3554] = -25;
        weight_rom[3555] = 1;
        weight_rom[3556] = -3;
        weight_rom[3557] = 3;
        weight_rom[3558] = -21;
        weight_rom[3559] = -16;
        weight_rom[3560] = -21;
        weight_rom[3561] = -37;
        weight_rom[3562] = -42;
        weight_rom[3563] = -23;
        weight_rom[3564] = -22;
        weight_rom[3565] = -5;
        weight_rom[3566] = -18;
        weight_rom[3567] = -4;
        weight_rom[3568] = 11;
        weight_rom[3569] = 28;
        weight_rom[3570] = 25;
        weight_rom[3571] = 19;
        weight_rom[3572] = 19;
        weight_rom[3573] = 7;
        weight_rom[3574] = -6;
        weight_rom[3575] = -26;
        weight_rom[3576] = -22;
        weight_rom[3577] = -39;
        weight_rom[3578] = -20;
        weight_rom[3579] = -15;
        weight_rom[3580] = -44;
        weight_rom[3581] = -31;
        weight_rom[3582] = -14;
        weight_rom[3583] = -4;
        weight_rom[3584] = 0;
        weight_rom[3585] = 3;
        weight_rom[3586] = -7;
        weight_rom[3587] = -15;
        weight_rom[3588] = -31;
        weight_rom[3589] = -50;
        weight_rom[3590] = -38;
        weight_rom[3591] = -18;
        weight_rom[3592] = -2;
        weight_rom[3593] = -3;
        weight_rom[3594] = 0;
        weight_rom[3595] = -4;
        weight_rom[3596] = 7;
        weight_rom[3597] = 15;
        weight_rom[3598] = 17;
        weight_rom[3599] = 8;
        weight_rom[3600] = 16;
        weight_rom[3601] = -10;
        weight_rom[3602] = -26;
        weight_rom[3603] = -37;
        weight_rom[3604] = -34;
        weight_rom[3605] = -37;
        weight_rom[3606] = -35;
        weight_rom[3607] = -22;
        weight_rom[3608] = -31;
        weight_rom[3609] = -43;
        weight_rom[3610] = -22;
        weight_rom[3611] = -2;
        weight_rom[3612] = 3;
        weight_rom[3613] = 14;
        weight_rom[3614] = -3;
        weight_rom[3615] = -27;
        weight_rom[3616] = -35;
        weight_rom[3617] = -46;
        weight_rom[3618] = -52;
        weight_rom[3619] = -10;
        weight_rom[3620] = 10;
        weight_rom[3621] = 7;
        weight_rom[3622] = -6;
        weight_rom[3623] = 0;
        weight_rom[3624] = 9;
        weight_rom[3625] = 9;
        weight_rom[3626] = 12;
        weight_rom[3627] = -9;
        weight_rom[3628] = -4;
        weight_rom[3629] = -20;
        weight_rom[3630] = -26;
        weight_rom[3631] = -23;
        weight_rom[3632] = -27;
        weight_rom[3633] = -13;
        weight_rom[3634] = -21;
        weight_rom[3635] = -17;
        weight_rom[3636] = -29;
        weight_rom[3637] = -53;
        weight_rom[3638] = -33;
        weight_rom[3639] = 0;
        weight_rom[3640] = 3;
        weight_rom[3641] = 11;
        weight_rom[3642] = -7;
        weight_rom[3643] = -33;
        weight_rom[3644] = -48;
        weight_rom[3645] = -45;
        weight_rom[3646] = -47;
        weight_rom[3647] = -26;
        weight_rom[3648] = -2;
        weight_rom[3649] = 4;
        weight_rom[3650] = -9;
        weight_rom[3651] = -5;
        weight_rom[3652] = -14;
        weight_rom[3653] = 0;
        weight_rom[3654] = -8;
        weight_rom[3655] = -13;
        weight_rom[3656] = -22;
        weight_rom[3657] = -19;
        weight_rom[3658] = -12;
        weight_rom[3659] = -15;
        weight_rom[3660] = -7;
        weight_rom[3661] = -18;
        weight_rom[3662] = -16;
        weight_rom[3663] = -23;
        weight_rom[3664] = -41;
        weight_rom[3665] = -31;
        weight_rom[3666] = 5;
        weight_rom[3667] = 8;
        weight_rom[3668] = 1;
        weight_rom[3669] = 7;
        weight_rom[3670] = -6;
        weight_rom[3671] = -27;
        weight_rom[3672] = -42;
        weight_rom[3673] = -32;
        weight_rom[3674] = -23;
        weight_rom[3675] = -19;
        weight_rom[3676] = -17;
        weight_rom[3677] = -7;
        weight_rom[3678] = -8;
        weight_rom[3679] = -23;
        weight_rom[3680] = -37;
        weight_rom[3681] = -26;
        weight_rom[3682] = -16;
        weight_rom[3683] = -20;
        weight_rom[3684] = -16;
        weight_rom[3685] = -20;
        weight_rom[3686] = -19;
        weight_rom[3687] = -13;
        weight_rom[3688] = -6;
        weight_rom[3689] = -18;
        weight_rom[3690] = -11;
        weight_rom[3691] = -7;
        weight_rom[3692] = -17;
        weight_rom[3693] = -20;
        weight_rom[3694] = -4;
        weight_rom[3695] = -3;
        weight_rom[3696] = 3;
        weight_rom[3697] = -5;
        weight_rom[3698] = -7;
        weight_rom[3699] = -28;
        weight_rom[3700] = -10;
        weight_rom[3701] = -13;
        weight_rom[3702] = -5;
        weight_rom[3703] = 6;
        weight_rom[3704] = -5;
        weight_rom[3705] = -10;
        weight_rom[3706] = -6;
        weight_rom[3707] = -23;
        weight_rom[3708] = -19;
        weight_rom[3709] = -14;
        weight_rom[3710] = -15;
        weight_rom[3711] = -9;
        weight_rom[3712] = -12;
        weight_rom[3713] = -10;
        weight_rom[3714] = -14;
        weight_rom[3715] = -14;
        weight_rom[3716] = -4;
        weight_rom[3717] = -1;
        weight_rom[3718] = -5;
        weight_rom[3719] = -11;
        weight_rom[3720] = -22;
        weight_rom[3721] = -8;
        weight_rom[3722] = -3;
        weight_rom[3723] = 1;
        weight_rom[3724] = 3;
        weight_rom[3725] = 7;
        weight_rom[3726] = -8;
        weight_rom[3727] = -47;
        weight_rom[3728] = -19;
        weight_rom[3729] = 3;
        weight_rom[3730] = 10;
        weight_rom[3731] = 3;
        weight_rom[3732] = -1;
        weight_rom[3733] = 6;
        weight_rom[3734] = 0;
        weight_rom[3735] = -6;
        weight_rom[3736] = -5;
        weight_rom[3737] = -12;
        weight_rom[3738] = -3;
        weight_rom[3739] = -5;
        weight_rom[3740] = -7;
        weight_rom[3741] = -15;
        weight_rom[3742] = -11;
        weight_rom[3743] = -9;
        weight_rom[3744] = -6;
        weight_rom[3745] = 6;
        weight_rom[3746] = -12;
        weight_rom[3747] = -31;
        weight_rom[3748] = -5;
        weight_rom[3749] = 5;
        weight_rom[3750] = -10;
        weight_rom[3751] = -1;
        weight_rom[3752] = 2;
        weight_rom[3753] = 0;
        weight_rom[3754] = -16;
        weight_rom[3755] = -22;
        weight_rom[3756] = -12;
        weight_rom[3757] = 15;
        weight_rom[3758] = 14;
        weight_rom[3759] = 15;
        weight_rom[3760] = 0;
        weight_rom[3761] = 1;
        weight_rom[3762] = 6;
        weight_rom[3763] = 6;
        weight_rom[3764] = 3;
        weight_rom[3765] = 9;
        weight_rom[3766] = 8;
        weight_rom[3767] = -2;
        weight_rom[3768] = 0;
        weight_rom[3769] = 3;
        weight_rom[3770] = -14;
        weight_rom[3771] = -14;
        weight_rom[3772] = -6;
        weight_rom[3773] = -11;
        weight_rom[3774] = -17;
        weight_rom[3775] = -6;
        weight_rom[3776] = -2;
        weight_rom[3777] = 11;
        weight_rom[3778] = 1;
        weight_rom[3779] = 4;
        weight_rom[3780] = -1;
        weight_rom[3781] = -3;
        weight_rom[3782] = -2;
        weight_rom[3783] = -19;
        weight_rom[3784] = -23;
        weight_rom[3785] = -14;
        weight_rom[3786] = -7;
        weight_rom[3787] = -1;
        weight_rom[3788] = 9;
        weight_rom[3789] = 0;
        weight_rom[3790] = -4;
        weight_rom[3791] = 3;
        weight_rom[3792] = 15;
        weight_rom[3793] = 19;
        weight_rom[3794] = 9;
        weight_rom[3795] = 5;
        weight_rom[3796] = 12;
        weight_rom[3797] = 14;
        weight_rom[3798] = -3;
        weight_rom[3799] = -6;
        weight_rom[3800] = -24;
        weight_rom[3801] = -12;
        weight_rom[3802] = -21;
        weight_rom[3803] = -8;
        weight_rom[3804] = -9;
        weight_rom[3805] = -11;
        weight_rom[3806] = 4;
        weight_rom[3807] = 2;
        weight_rom[3808] = 4;
        weight_rom[3809] = -3;
        weight_rom[3810] = -9;
        weight_rom[3811] = -35;
        weight_rom[3812] = -34;
        weight_rom[3813] = -4;
        weight_rom[3814] = -10;
        weight_rom[3815] = 0;
        weight_rom[3816] = 5;
        weight_rom[3817] = -1;
        weight_rom[3818] = 6;
        weight_rom[3819] = 4;
        weight_rom[3820] = 0;
        weight_rom[3821] = -14;
        weight_rom[3822] = -13;
        weight_rom[3823] = 5;
        weight_rom[3824] = 9;
        weight_rom[3825] = -8;
        weight_rom[3826] = 14;
        weight_rom[3827] = 13;
        weight_rom[3828] = -3;
        weight_rom[3829] = -17;
        weight_rom[3830] = -11;
        weight_rom[3831] = 2;
        weight_rom[3832] = -16;
        weight_rom[3833] = -26;
        weight_rom[3834] = 2;
        weight_rom[3835] = 2;
        weight_rom[3836] = 0;
        weight_rom[3837] = -1;
        weight_rom[3838] = -4;
        weight_rom[3839] = 1;
        weight_rom[3840] = -8;
        weight_rom[3841] = -5;
        weight_rom[3842] = -19;
        weight_rom[3843] = -1;
        weight_rom[3844] = -11;
        weight_rom[3845] = -9;
        weight_rom[3846] = -15;
        weight_rom[3847] = -10;
        weight_rom[3848] = -23;
        weight_rom[3849] = -5;
        weight_rom[3850] = 0;
        weight_rom[3851] = -5;
        weight_rom[3852] = 3;
        weight_rom[3853] = 1;
        weight_rom[3854] = 11;
        weight_rom[3855] = 6;
        weight_rom[3856] = 5;
        weight_rom[3857] = -6;
        weight_rom[3858] = -14;
        weight_rom[3859] = -9;
        weight_rom[3860] = 3;
        weight_rom[3861] = -2;
        weight_rom[3862] = 2;
        weight_rom[3863] = -3;
        weight_rom[3864] = -3;
        weight_rom[3865] = -1;
        weight_rom[3866] = 3;
        weight_rom[3867] = 0;
        weight_rom[3868] = 20;
        weight_rom[3869] = 33;
        weight_rom[3870] = 20;
        weight_rom[3871] = 22;
        weight_rom[3872] = 22;
        weight_rom[3873] = 12;
        weight_rom[3874] = 3;
        weight_rom[3875] = -1;
        weight_rom[3876] = -2;
        weight_rom[3877] = 4;
        weight_rom[3878] = 13;
        weight_rom[3879] = -1;
        weight_rom[3880] = 5;
        weight_rom[3881] = 15;
        weight_rom[3882] = 20;
        weight_rom[3883] = 4;
        weight_rom[3884] = 4;
        weight_rom[3885] = 1;
        weight_rom[3886] = -2;
        weight_rom[3887] = 6;
        weight_rom[3888] = 0;
        weight_rom[3889] = -2;
        weight_rom[3890] = 2;
        weight_rom[3891] = -2;
        weight_rom[3892] = 3;
        weight_rom[3893] = -1;
        weight_rom[3894] = -3;
        weight_rom[3895] = 3;
        weight_rom[3896] = -4;
        weight_rom[3897] = -18;
        weight_rom[3898] = -33;
        weight_rom[3899] = 6;
        weight_rom[3900] = 1;
        weight_rom[3901] = -2;
        weight_rom[3902] = -6;
        weight_rom[3903] = 3;
        weight_rom[3904] = 4;
        weight_rom[3905] = -29;
        weight_rom[3906] = 1;
        weight_rom[3907] = 8;
        weight_rom[3908] = 2;
        weight_rom[3909] = -28;
        weight_rom[3910] = -3;
        weight_rom[3911] = 6;
        weight_rom[3912] = -6;
        weight_rom[3913] = -7;
        weight_rom[3914] = 0;
        weight_rom[3915] = 0;
        weight_rom[3916] = 3;
        weight_rom[3917] = 3;
        weight_rom[3918] = -1;
        weight_rom[3919] = 3;
        weight_rom[3920] = -4;
        weight_rom[3921] = 2;
        weight_rom[3922] = 4;
        weight_rom[3923] = -1;
        weight_rom[3924] = -2;
        weight_rom[3925] = -1;
        weight_rom[3926] = 0;
        weight_rom[3927] = 4;
        weight_rom[3928] = 3;
        weight_rom[3929] = 4;
        weight_rom[3930] = 2;
        weight_rom[3931] = 4;
        weight_rom[3932] = -3;
        weight_rom[3933] = -11;
        weight_rom[3934] = 2;
        weight_rom[3935] = 4;
        weight_rom[3936] = 1;
        weight_rom[3937] = -2;
        weight_rom[3938] = 2;
        weight_rom[3939] = -4;
        weight_rom[3940] = 3;
        weight_rom[3941] = 4;
        weight_rom[3942] = -2;
        weight_rom[3943] = -4;
        weight_rom[3944] = 1;
        weight_rom[3945] = 4;
        weight_rom[3946] = -3;
        weight_rom[3947] = 0;
        weight_rom[3948] = 3;
        weight_rom[3949] = 2;
        weight_rom[3950] = -3;
        weight_rom[3951] = -4;
        weight_rom[3952] = 0;
        weight_rom[3953] = 0;
        weight_rom[3954] = -14;
        weight_rom[3955] = -28;
        weight_rom[3956] = -21;
        weight_rom[3957] = -11;
        weight_rom[3958] = -20;
        weight_rom[3959] = -16;
        weight_rom[3960] = -34;
        weight_rom[3961] = -24;
        weight_rom[3962] = 1;
        weight_rom[3963] = -24;
        weight_rom[3964] = -36;
        weight_rom[3965] = -32;
        weight_rom[3966] = -26;
        weight_rom[3967] = -22;
        weight_rom[3968] = -22;
        weight_rom[3969] = -17;
        weight_rom[3970] = -18;
        weight_rom[3971] = -12;
        weight_rom[3972] = 1;
        weight_rom[3973] = 0;
        weight_rom[3974] = -3;
        weight_rom[3975] = 4;
        weight_rom[3976] = -3;
        weight_rom[3977] = -4;
        weight_rom[3978] = 2;
        weight_rom[3979] = 0;
        weight_rom[3980] = -18;
        weight_rom[3981] = 1;
        weight_rom[3982] = -29;
        weight_rom[3983] = -44;
        weight_rom[3984] = -38;
        weight_rom[3985] = -52;
        weight_rom[3986] = -60;
        weight_rom[3987] = -63;
        weight_rom[3988] = -67;
        weight_rom[3989] = -53;
        weight_rom[3990] = -62;
        weight_rom[3991] = -51;
        weight_rom[3992] = -25;
        weight_rom[3993] = -28;
        weight_rom[3994] = -3;
        weight_rom[3995] = 1;
        weight_rom[3996] = -17;
        weight_rom[3997] = -19;
        weight_rom[3998] = -22;
        weight_rom[3999] = -25;
        weight_rom[4000] = -28;
        weight_rom[4001] = -19;
        weight_rom[4002] = -2;
        weight_rom[4003] = 3;
        weight_rom[4004] = 0;
        weight_rom[4005] = 2;
        weight_rom[4006] = -6;
        weight_rom[4007] = 3;
        weight_rom[4008] = 5;
        weight_rom[4009] = -4;
        weight_rom[4010] = -32;
        weight_rom[4011] = -20;
        weight_rom[4012] = -36;
        weight_rom[4013] = -58;
        weight_rom[4014] = -42;
        weight_rom[4015] = -62;
        weight_rom[4016] = -46;
        weight_rom[4017] = -39;
        weight_rom[4018] = -18;
        weight_rom[4019] = -28;
        weight_rom[4020] = -20;
        weight_rom[4021] = -13;
        weight_rom[4022] = -15;
        weight_rom[4023] = -9;
        weight_rom[4024] = 7;
        weight_rom[4025] = 7;
        weight_rom[4026] = 12;
        weight_rom[4027] = -6;
        weight_rom[4028] = -12;
        weight_rom[4029] = 16;
        weight_rom[4030] = -2;
        weight_rom[4031] = -3;
        weight_rom[4032] = -3;
        weight_rom[4033] = -1;
        weight_rom[4034] = 8;
        weight_rom[4035] = -4;
        weight_rom[4036] = -3;
        weight_rom[4037] = -16;
        weight_rom[4038] = -11;
        weight_rom[4039] = -9;
        weight_rom[4040] = -16;
        weight_rom[4041] = -9;
        weight_rom[4042] = -19;
        weight_rom[4043] = 3;
        weight_rom[4044] = 2;
        weight_rom[4045] = -13;
        weight_rom[4046] = 2;
        weight_rom[4047] = -1;
        weight_rom[4048] = 7;
        weight_rom[4049] = -5;
        weight_rom[4050] = -2;
        weight_rom[4051] = -5;
        weight_rom[4052] = -3;
        weight_rom[4053] = 23;
        weight_rom[4054] = 6;
        weight_rom[4055] = 15;
        weight_rom[4056] = 35;
        weight_rom[4057] = 19;
        weight_rom[4058] = 14;
        weight_rom[4059] = -1;
        weight_rom[4060] = 4;
        weight_rom[4061] = -3;
        weight_rom[4062] = -1;
        weight_rom[4063] = 5;
        weight_rom[4064] = -26;
        weight_rom[4065] = 7;
        weight_rom[4066] = -2;
        weight_rom[4067] = 7;
        weight_rom[4068] = 16;
        weight_rom[4069] = 24;
        weight_rom[4070] = 12;
        weight_rom[4071] = 19;
        weight_rom[4072] = 13;
        weight_rom[4073] = 4;
        weight_rom[4074] = -5;
        weight_rom[4075] = -2;
        weight_rom[4076] = 2;
        weight_rom[4077] = -1;
        weight_rom[4078] = -22;
        weight_rom[4079] = -18;
        weight_rom[4080] = -5;
        weight_rom[4081] = 2;
        weight_rom[4082] = 1;
        weight_rom[4083] = 13;
        weight_rom[4084] = 3;
        weight_rom[4085] = 32;
        weight_rom[4086] = 0;
        weight_rom[4087] = 2;
        weight_rom[4088] = 0;
        weight_rom[4089] = 3;
        weight_rom[4090] = 13;
        weight_rom[4091] = -5;
        weight_rom[4092] = 10;
        weight_rom[4093] = 10;
        weight_rom[4094] = 19;
        weight_rom[4095] = 14;
        weight_rom[4096] = 26;
        weight_rom[4097] = 21;
        weight_rom[4098] = 16;
        weight_rom[4099] = 13;
        weight_rom[4100] = 11;
        weight_rom[4101] = -5;
        weight_rom[4102] = -11;
        weight_rom[4103] = 5;
        weight_rom[4104] = -10;
        weight_rom[4105] = -7;
        weight_rom[4106] = -25;
        weight_rom[4107] = -4;
        weight_rom[4108] = -3;
        weight_rom[4109] = 9;
        weight_rom[4110] = 7;
        weight_rom[4111] = 15;
        weight_rom[4112] = 42;
        weight_rom[4113] = 40;
        weight_rom[4114] = 18;
        weight_rom[4115] = -5;
        weight_rom[4116] = 2;
        weight_rom[4117] = -11;
        weight_rom[4118] = 8;
        weight_rom[4119] = 8;
        weight_rom[4120] = -10;
        weight_rom[4121] = 9;
        weight_rom[4122] = 11;
        weight_rom[4123] = 28;
        weight_rom[4124] = 24;
        weight_rom[4125] = 15;
        weight_rom[4126] = 17;
        weight_rom[4127] = 12;
        weight_rom[4128] = 4;
        weight_rom[4129] = -3;
        weight_rom[4130] = -16;
        weight_rom[4131] = -4;
        weight_rom[4132] = 0;
        weight_rom[4133] = 3;
        weight_rom[4134] = -1;
        weight_rom[4135] = -1;
        weight_rom[4136] = 4;
        weight_rom[4137] = 11;
        weight_rom[4138] = 13;
        weight_rom[4139] = 39;
        weight_rom[4140] = 37;
        weight_rom[4141] = 43;
        weight_rom[4142] = 8;
        weight_rom[4143] = 8;
        weight_rom[4144] = 14;
        weight_rom[4145] = 12;
        weight_rom[4146] = 4;
        weight_rom[4147] = 12;
        weight_rom[4148] = -2;
        weight_rom[4149] = 10;
        weight_rom[4150] = 20;
        weight_rom[4151] = 28;
        weight_rom[4152] = 17;
        weight_rom[4153] = 17;
        weight_rom[4154] = 13;
        weight_rom[4155] = 9;
        weight_rom[4156] = 15;
        weight_rom[4157] = 6;
        weight_rom[4158] = -5;
        weight_rom[4159] = 4;
        weight_rom[4160] = 14;
        weight_rom[4161] = -2;
        weight_rom[4162] = 9;
        weight_rom[4163] = -2;
        weight_rom[4164] = 11;
        weight_rom[4165] = 9;
        weight_rom[4166] = 21;
        weight_rom[4167] = 47;
        weight_rom[4168] = 71;
        weight_rom[4169] = 64;
        weight_rom[4170] = 45;
        weight_rom[4171] = 11;
        weight_rom[4172] = 12;
        weight_rom[4173] = 12;
        weight_rom[4174] = 10;
        weight_rom[4175] = 6;
        weight_rom[4176] = -5;
        weight_rom[4177] = 11;
        weight_rom[4178] = 8;
        weight_rom[4179] = 9;
        weight_rom[4180] = 22;
        weight_rom[4181] = 21;
        weight_rom[4182] = 17;
        weight_rom[4183] = 23;
        weight_rom[4184] = 20;
        weight_rom[4185] = 10;
        weight_rom[4186] = 8;
        weight_rom[4187] = -4;
        weight_rom[4188] = 2;
        weight_rom[4189] = 1;
        weight_rom[4190] = 1;
        weight_rom[4191] = 3;
        weight_rom[4192] = 13;
        weight_rom[4193] = 22;
        weight_rom[4194] = 25;
        weight_rom[4195] = 32;
        weight_rom[4196] = 60;
        weight_rom[4197] = 81;
        weight_rom[4198] = 41;
        weight_rom[4199] = 17;
        weight_rom[4200] = 17;
        weight_rom[4201] = 20;
        weight_rom[4202] = 22;
        weight_rom[4203] = 1;
        weight_rom[4204] = 11;
        weight_rom[4205] = -8;
        weight_rom[4206] = 3;
        weight_rom[4207] = 19;
        weight_rom[4208] = 19;
        weight_rom[4209] = 30;
        weight_rom[4210] = 21;
        weight_rom[4211] = 22;
        weight_rom[4212] = 23;
        weight_rom[4213] = 22;
        weight_rom[4214] = 18;
        weight_rom[4215] = 10;
        weight_rom[4216] = 6;
        weight_rom[4217] = -7;
        weight_rom[4218] = -2;
        weight_rom[4219] = 16;
        weight_rom[4220] = 14;
        weight_rom[4221] = 27;
        weight_rom[4222] = 18;
        weight_rom[4223] = 36;
        weight_rom[4224] = 50;
        weight_rom[4225] = 73;
        weight_rom[4226] = 51;
        weight_rom[4227] = 15;
        weight_rom[4228] = 21;
        weight_rom[4229] = 20;
        weight_rom[4230] = 31;
        weight_rom[4231] = -6;
        weight_rom[4232] = 11;
        weight_rom[4233] = 2;
        weight_rom[4234] = 23;
        weight_rom[4235] = 19;
        weight_rom[4236] = 20;
        weight_rom[4237] = 26;
        weight_rom[4238] = 26;
        weight_rom[4239] = 24;
        weight_rom[4240] = 32;
        weight_rom[4241] = 26;
        weight_rom[4242] = 27;
        weight_rom[4243] = 24;
        weight_rom[4244] = 11;
        weight_rom[4245] = 3;
        weight_rom[4246] = 6;
        weight_rom[4247] = -3;
        weight_rom[4248] = -1;
        weight_rom[4249] = -3;
        weight_rom[4250] = 17;
        weight_rom[4251] = 18;
        weight_rom[4252] = 26;
        weight_rom[4253] = 48;
        weight_rom[4254] = 57;
        weight_rom[4255] = 2;
        weight_rom[4256] = 16;
        weight_rom[4257] = 15;
        weight_rom[4258] = 22;
        weight_rom[4259] = 20;
        weight_rom[4260] = 11;
        weight_rom[4261] = 6;
        weight_rom[4262] = 7;
        weight_rom[4263] = 20;
        weight_rom[4264] = 26;
        weight_rom[4265] = 19;
        weight_rom[4266] = 23;
        weight_rom[4267] = 26;
        weight_rom[4268] = 19;
        weight_rom[4269] = 14;
        weight_rom[4270] = 13;
        weight_rom[4271] = 21;
        weight_rom[4272] = 4;
        weight_rom[4273] = 2;
        weight_rom[4274] = 1;
        weight_rom[4275] = 0;
        weight_rom[4276] = 10;
        weight_rom[4277] = 0;
        weight_rom[4278] = -18;
        weight_rom[4279] = -22;
        weight_rom[4280] = -32;
        weight_rom[4281] = 11;
        weight_rom[4282] = 37;
        weight_rom[4283] = -3;
        weight_rom[4284] = 1;
        weight_rom[4285] = 9;
        weight_rom[4286] = 32;
        weight_rom[4287] = 8;
        weight_rom[4288] = 11;
        weight_rom[4289] = 0;
        weight_rom[4290] = -3;
        weight_rom[4291] = 2;
        weight_rom[4292] = 0;
        weight_rom[4293] = 4;
        weight_rom[4294] = 17;
        weight_rom[4295] = 24;
        weight_rom[4296] = 19;
        weight_rom[4297] = 12;
        weight_rom[4298] = -7;
        weight_rom[4299] = 8;
        weight_rom[4300] = 0;
        weight_rom[4301] = -5;
        weight_rom[4302] = 8;
        weight_rom[4303] = 8;
        weight_rom[4304] = 10;
        weight_rom[4305] = 0;
        weight_rom[4306] = -4;
        weight_rom[4307] = -27;
        weight_rom[4308] = -18;
        weight_rom[4309] = -11;
        weight_rom[4310] = 1;
        weight_rom[4311] = -24;
        weight_rom[4312] = 3;
        weight_rom[4313] = 10;
        weight_rom[4314] = 19;
        weight_rom[4315] = 2;
        weight_rom[4316] = 4;
        weight_rom[4317] = -10;
        weight_rom[4318] = -20;
        weight_rom[4319] = -23;
        weight_rom[4320] = -19;
        weight_rom[4321] = -12;
        weight_rom[4322] = 15;
        weight_rom[4323] = 10;
        weight_rom[4324] = 10;
        weight_rom[4325] = 13;
        weight_rom[4326] = 6;
        weight_rom[4327] = -3;
        weight_rom[4328] = 2;
        weight_rom[4329] = 11;
        weight_rom[4330] = 3;
        weight_rom[4331] = 13;
        weight_rom[4332] = 6;
        weight_rom[4333] = -8;
        weight_rom[4334] = 6;
        weight_rom[4335] = 0;
        weight_rom[4336] = -12;
        weight_rom[4337] = -19;
        weight_rom[4338] = -33;
        weight_rom[4339] = -4;
        weight_rom[4340] = 4;
        weight_rom[4341] = 6;
        weight_rom[4342] = 25;
        weight_rom[4343] = 1;
        weight_rom[4344] = -18;
        weight_rom[4345] = -26;
        weight_rom[4346] = -13;
        weight_rom[4347] = -35;
        weight_rom[4348] = -25;
        weight_rom[4349] = -14;
        weight_rom[4350] = -2;
        weight_rom[4351] = -3;
        weight_rom[4352] = 7;
        weight_rom[4353] = 2;
        weight_rom[4354] = 0;
        weight_rom[4355] = 6;
        weight_rom[4356] = 10;
        weight_rom[4357] = 19;
        weight_rom[4358] = 16;
        weight_rom[4359] = 1;
        weight_rom[4360] = 3;
        weight_rom[4361] = 9;
        weight_rom[4362] = 13;
        weight_rom[4363] = 11;
        weight_rom[4364] = -7;
        weight_rom[4365] = -35;
        weight_rom[4366] = -19;
        weight_rom[4367] = -13;
        weight_rom[4368] = -4;
        weight_rom[4369] = 1;
        weight_rom[4370] = -13;
        weight_rom[4371] = -3;
        weight_rom[4372] = -18;
        weight_rom[4373] = -33;
        weight_rom[4374] = -9;
        weight_rom[4375] = -24;
        weight_rom[4376] = -14;
        weight_rom[4377] = -25;
        weight_rom[4378] = -32;
        weight_rom[4379] = -27;
        weight_rom[4380] = 1;
        weight_rom[4381] = 3;
        weight_rom[4382] = 0;
        weight_rom[4383] = 15;
        weight_rom[4384] = 18;
        weight_rom[4385] = 11;
        weight_rom[4386] = -4;
        weight_rom[4387] = -13;
        weight_rom[4388] = -11;
        weight_rom[4389] = -3;
        weight_rom[4390] = 10;
        weight_rom[4391] = 12;
        weight_rom[4392] = -4;
        weight_rom[4393] = -33;
        weight_rom[4394] = -26;
        weight_rom[4395] = -12;
        weight_rom[4396] = 2;
        weight_rom[4397] = 4;
        weight_rom[4398] = -22;
        weight_rom[4399] = -15;
        weight_rom[4400] = 2;
        weight_rom[4401] = -2;
        weight_rom[4402] = 6;
        weight_rom[4403] = -9;
        weight_rom[4404] = -11;
        weight_rom[4405] = -7;
        weight_rom[4406] = -22;
        weight_rom[4407] = -17;
        weight_rom[4408] = -7;
        weight_rom[4409] = 1;
        weight_rom[4410] = 17;
        weight_rom[4411] = 14;
        weight_rom[4412] = 13;
        weight_rom[4413] = 1;
        weight_rom[4414] = -7;
        weight_rom[4415] = -15;
        weight_rom[4416] = -5;
        weight_rom[4417] = 10;
        weight_rom[4418] = 1;
        weight_rom[4419] = 9;
        weight_rom[4420] = 19;
        weight_rom[4421] = -38;
        weight_rom[4422] = -31;
        weight_rom[4423] = 2;
        weight_rom[4424] = -3;
        weight_rom[4425] = -3;
        weight_rom[4426] = -3;
        weight_rom[4427] = -8;
        weight_rom[4428] = 7;
        weight_rom[4429] = 13;
        weight_rom[4430] = 10;
        weight_rom[4431] = -13;
        weight_rom[4432] = -6;
        weight_rom[4433] = -11;
        weight_rom[4434] = -15;
        weight_rom[4435] = -1;
        weight_rom[4436] = -11;
        weight_rom[4437] = 12;
        weight_rom[4438] = 17;
        weight_rom[4439] = 12;
        weight_rom[4440] = -10;
        weight_rom[4441] = -17;
        weight_rom[4442] = -22;
        weight_rom[4443] = -15;
        weight_rom[4444] = -4;
        weight_rom[4445] = -6;
        weight_rom[4446] = 1;
        weight_rom[4447] = 1;
        weight_rom[4448] = -7;
        weight_rom[4449] = -48;
        weight_rom[4450] = -20;
        weight_rom[4451] = -10;
        weight_rom[4452] = -3;
        weight_rom[4453] = 0;
        weight_rom[4454] = -3;
        weight_rom[4455] = -11;
        weight_rom[4456] = 10;
        weight_rom[4457] = 24;
        weight_rom[4458] = -2;
        weight_rom[4459] = -11;
        weight_rom[4460] = -1;
        weight_rom[4461] = -8;
        weight_rom[4462] = -15;
        weight_rom[4463] = -20;
        weight_rom[4464] = -2;
        weight_rom[4465] = -3;
        weight_rom[4466] = 5;
        weight_rom[4467] = -9;
        weight_rom[4468] = -24;
        weight_rom[4469] = -27;
        weight_rom[4470] = -24;
        weight_rom[4471] = -18;
        weight_rom[4472] = -14;
        weight_rom[4473] = -11;
        weight_rom[4474] = -4;
        weight_rom[4475] = 14;
        weight_rom[4476] = 25;
        weight_rom[4477] = 0;
        weight_rom[4478] = -24;
        weight_rom[4479] = 4;
        weight_rom[4480] = 3;
        weight_rom[4481] = -22;
        weight_rom[4482] = -19;
        weight_rom[4483] = -21;
        weight_rom[4484] = -25;
        weight_rom[4485] = 5;
        weight_rom[4486] = 0;
        weight_rom[4487] = -10;
        weight_rom[4488] = -12;
        weight_rom[4489] = -17;
        weight_rom[4490] = -18;
        weight_rom[4491] = -11;
        weight_rom[4492] = -6;
        weight_rom[4493] = 4;
        weight_rom[4494] = -5;
        weight_rom[4495] = -8;
        weight_rom[4496] = -20;
        weight_rom[4497] = -17;
        weight_rom[4498] = -32;
        weight_rom[4499] = -17;
        weight_rom[4500] = -15;
        weight_rom[4501] = -9;
        weight_rom[4502] = 6;
        weight_rom[4503] = 15;
        weight_rom[4504] = 4;
        weight_rom[4505] = 0;
        weight_rom[4506] = -21;
        weight_rom[4507] = -1;
        weight_rom[4508] = -1;
        weight_rom[4509] = -13;
        weight_rom[4510] = -19;
        weight_rom[4511] = -36;
        weight_rom[4512] = -14;
        weight_rom[4513] = -4;
        weight_rom[4514] = 10;
        weight_rom[4515] = -2;
        weight_rom[4516] = 1;
        weight_rom[4517] = 0;
        weight_rom[4518] = -13;
        weight_rom[4519] = -7;
        weight_rom[4520] = -2;
        weight_rom[4521] = -4;
        weight_rom[4522] = -8;
        weight_rom[4523] = 0;
        weight_rom[4524] = -15;
        weight_rom[4525] = -16;
        weight_rom[4526] = -24;
        weight_rom[4527] = -19;
        weight_rom[4528] = -8;
        weight_rom[4529] = -1;
        weight_rom[4530] = 8;
        weight_rom[4531] = -3;
        weight_rom[4532] = -13;
        weight_rom[4533] = -5;
        weight_rom[4534] = -17;
        weight_rom[4535] = -4;
        weight_rom[4536] = 2;
        weight_rom[4537] = 5;
        weight_rom[4538] = -14;
        weight_rom[4539] = -42;
        weight_rom[4540] = -8;
        weight_rom[4541] = -7;
        weight_rom[4542] = -5;
        weight_rom[4543] = 17;
        weight_rom[4544] = 0;
        weight_rom[4545] = 0;
        weight_rom[4546] = 2;
        weight_rom[4547] = 5;
        weight_rom[4548] = 5;
        weight_rom[4549] = 7;
        weight_rom[4550] = 0;
        weight_rom[4551] = -5;
        weight_rom[4552] = -7;
        weight_rom[4553] = -10;
        weight_rom[4554] = -15;
        weight_rom[4555] = -14;
        weight_rom[4556] = -19;
        weight_rom[4557] = -6;
        weight_rom[4558] = -10;
        weight_rom[4559] = 1;
        weight_rom[4560] = 2;
        weight_rom[4561] = 3;
        weight_rom[4562] = -3;
        weight_rom[4563] = -4;
        weight_rom[4564] = 2;
        weight_rom[4565] = -3;
        weight_rom[4566] = -14;
        weight_rom[4567] = -18;
        weight_rom[4568] = 7;
        weight_rom[4569] = 6;
        weight_rom[4570] = 2;
        weight_rom[4571] = 11;
        weight_rom[4572] = -4;
        weight_rom[4573] = 16;
        weight_rom[4574] = 15;
        weight_rom[4575] = 13;
        weight_rom[4576] = 12;
        weight_rom[4577] = 8;
        weight_rom[4578] = 11;
        weight_rom[4579] = 11;
        weight_rom[4580] = 9;
        weight_rom[4581] = -4;
        weight_rom[4582] = -20;
        weight_rom[4583] = -11;
        weight_rom[4584] = -21;
        weight_rom[4585] = -19;
        weight_rom[4586] = -15;
        weight_rom[4587] = -8;
        weight_rom[4588] = 5;
        weight_rom[4589] = 3;
        weight_rom[4590] = -12;
        weight_rom[4591] = -4;
        weight_rom[4592] = 4;
        weight_rom[4593] = -2;
        weight_rom[4594] = -7;
        weight_rom[4595] = 20;
        weight_rom[4596] = -12;
        weight_rom[4597] = 19;
        weight_rom[4598] = 4;
        weight_rom[4599] = 14;
        weight_rom[4600] = 26;
        weight_rom[4601] = 16;
        weight_rom[4602] = 18;
        weight_rom[4603] = 30;
        weight_rom[4604] = 26;
        weight_rom[4605] = 29;
        weight_rom[4606] = 22;
        weight_rom[4607] = 22;
        weight_rom[4608] = 14;
        weight_rom[4609] = -7;
        weight_rom[4610] = -3;
        weight_rom[4611] = 0;
        weight_rom[4612] = -14;
        weight_rom[4613] = -18;
        weight_rom[4614] = -22;
        weight_rom[4615] = -2;
        weight_rom[4616] = -11;
        weight_rom[4617] = -26;
        weight_rom[4618] = 3;
        weight_rom[4619] = 0;
        weight_rom[4620] = -3;
        weight_rom[4621] = 3;
        weight_rom[4622] = 2;
        weight_rom[4623] = 20;
        weight_rom[4624] = 17;
        weight_rom[4625] = -3;
        weight_rom[4626] = 7;
        weight_rom[4627] = 9;
        weight_rom[4628] = 12;
        weight_rom[4629] = 21;
        weight_rom[4630] = 27;
        weight_rom[4631] = 33;
        weight_rom[4632] = 26;
        weight_rom[4633] = 26;
        weight_rom[4634] = 28;
        weight_rom[4635] = 37;
        weight_rom[4636] = 23;
        weight_rom[4637] = 19;
        weight_rom[4638] = 15;
        weight_rom[4639] = 3;
        weight_rom[4640] = -14;
        weight_rom[4641] = 0;
        weight_rom[4642] = 9;
        weight_rom[4643] = 14;
        weight_rom[4644] = 9;
        weight_rom[4645] = 1;
        weight_rom[4646] = 1;
        weight_rom[4647] = -4;
        weight_rom[4648] = -4;
        weight_rom[4649] = 3;
        weight_rom[4650] = -1;
        weight_rom[4651] = -4;
        weight_rom[4652] = -27;
        weight_rom[4653] = -21;
        weight_rom[4654] = -16;
        weight_rom[4655] = -7;
        weight_rom[4656] = -1;
        weight_rom[4657] = 12;
        weight_rom[4658] = 9;
        weight_rom[4659] = 20;
        weight_rom[4660] = 7;
        weight_rom[4661] = 23;
        weight_rom[4662] = 9;
        weight_rom[4663] = 23;
        weight_rom[4664] = 17;
        weight_rom[4665] = 16;
        weight_rom[4666] = 1;
        weight_rom[4667] = 12;
        weight_rom[4668] = -1;
        weight_rom[4669] = -3;
        weight_rom[4670] = 14;
        weight_rom[4671] = -8;
        weight_rom[4672] = 0;
        weight_rom[4673] = -2;
        weight_rom[4674] = 2;
        weight_rom[4675] = -2;
        weight_rom[4676] = -1;
        weight_rom[4677] = 1;
        weight_rom[4678] = 1;
        weight_rom[4679] = 2;
        weight_rom[4680] = 4;
        weight_rom[4681] = 25;
        weight_rom[4682] = 20;
        weight_rom[4683] = -5;
        weight_rom[4684] = 5;
        weight_rom[4685] = 5;
        weight_rom[4686] = 19;
        weight_rom[4687] = 9;
        weight_rom[4688] = 4;
        weight_rom[4689] = 36;
        weight_rom[4690] = 16;
        weight_rom[4691] = 5;
        weight_rom[4692] = 8;
        weight_rom[4693] = 38;
        weight_rom[4694] = 20;
        weight_rom[4695] = -3;
        weight_rom[4696] = 6;
        weight_rom[4697] = 3;
        weight_rom[4698] = 9;
        weight_rom[4699] = -1;
        weight_rom[4700] = -1;
        weight_rom[4701] = 1;
        weight_rom[4702] = 1;
        weight_rom[4703] = 4;
        weight_rom[4704] = 1;
        weight_rom[4705] = 4;
        weight_rom[4706] = 2;
        weight_rom[4707] = -2;
        weight_rom[4708] = 0;
        weight_rom[4709] = -2;
        weight_rom[4710] = -3;
        weight_rom[4711] = 3;
        weight_rom[4712] = 1;
        weight_rom[4713] = -2;
        weight_rom[4714] = 5;
        weight_rom[4715] = -1;
        weight_rom[4716] = 2;
        weight_rom[4717] = 4;
        weight_rom[4718] = 9;
        weight_rom[4719] = -3;
        weight_rom[4720] = -2;
        weight_rom[4721] = 2;
        weight_rom[4722] = 4;
        weight_rom[4723] = -3;
        weight_rom[4724] = -4;
        weight_rom[4725] = -2;
        weight_rom[4726] = -3;
        weight_rom[4727] = 3;
        weight_rom[4728] = -2;
        weight_rom[4729] = 0;
        weight_rom[4730] = 2;
        weight_rom[4731] = 0;
        weight_rom[4732] = 1;
        weight_rom[4733] = 3;
        weight_rom[4734] = 4;
        weight_rom[4735] = -2;
        weight_rom[4736] = -4;
        weight_rom[4737] = -4;
        weight_rom[4738] = 5;
        weight_rom[4739] = 1;
        weight_rom[4740] = 2;
        weight_rom[4741] = -5;
        weight_rom[4742] = -6;
        weight_rom[4743] = 10;
        weight_rom[4744] = 6;
        weight_rom[4745] = -13;
        weight_rom[4746] = 4;
        weight_rom[4747] = 10;
        weight_rom[4748] = 32;
        weight_rom[4749] = -7;
        weight_rom[4750] = -14;
        weight_rom[4751] = -15;
        weight_rom[4752] = -7;
        weight_rom[4753] = -3;
        weight_rom[4754] = -3;
        weight_rom[4755] = -4;
        weight_rom[4756] = 2;
        weight_rom[4757] = 4;
        weight_rom[4758] = 2;
        weight_rom[4759] = 4;
        weight_rom[4760] = 3;
        weight_rom[4761] = 4;
        weight_rom[4762] = -3;
        weight_rom[4763] = -3;
        weight_rom[4764] = -1;
        weight_rom[4765] = 3;
        weight_rom[4766] = -9;
        weight_rom[4767] = -7;
        weight_rom[4768] = -10;
        weight_rom[4769] = -3;
        weight_rom[4770] = -19;
        weight_rom[4771] = -9;
        weight_rom[4772] = -5;
        weight_rom[4773] = 7;
        weight_rom[4774] = -5;
        weight_rom[4775] = -13;
        weight_rom[4776] = 8;
        weight_rom[4777] = -14;
        weight_rom[4778] = -32;
        weight_rom[4779] = -36;
        weight_rom[4780] = -17;
        weight_rom[4781] = -15;
        weight_rom[4782] = -24;
        weight_rom[4783] = -4;
        weight_rom[4784] = 8;
        weight_rom[4785] = 10;
        weight_rom[4786] = 2;
        weight_rom[4787] = 1;
        weight_rom[4788] = -4;
        weight_rom[4789] = 0;
        weight_rom[4790] = -5;
        weight_rom[4791] = 1;
        weight_rom[4792] = 1;
        weight_rom[4793] = 14;
        weight_rom[4794] = -14;
        weight_rom[4795] = -2;
        weight_rom[4796] = 13;
        weight_rom[4797] = -1;
        weight_rom[4798] = 3;
        weight_rom[4799] = 28;
        weight_rom[4800] = 43;
        weight_rom[4801] = 34;
        weight_rom[4802] = 36;
        weight_rom[4803] = 5;
        weight_rom[4804] = 6;
        weight_rom[4805] = 6;
        weight_rom[4806] = -17;
        weight_rom[4807] = -35;
        weight_rom[4808] = -25;
        weight_rom[4809] = -53;
        weight_rom[4810] = -37;
        weight_rom[4811] = -28;
        weight_rom[4812] = -11;
        weight_rom[4813] = 16;
        weight_rom[4814] = -1;
        weight_rom[4815] = 1;
        weight_rom[4816] = 0;
        weight_rom[4817] = 0;
        weight_rom[4818] = 9;
        weight_rom[4819] = -2;
        weight_rom[4820] = -10;
        weight_rom[4821] = 5;
        weight_rom[4822] = 22;
        weight_rom[4823] = -5;
        weight_rom[4824] = 3;
        weight_rom[4825] = 16;
        weight_rom[4826] = 20;
        weight_rom[4827] = 28;
        weight_rom[4828] = 30;
        weight_rom[4829] = 27;
        weight_rom[4830] = 33;
        weight_rom[4831] = 28;
        weight_rom[4832] = 10;
        weight_rom[4833] = 5;
        weight_rom[4834] = 12;
        weight_rom[4835] = -13;
        weight_rom[4836] = -15;
        weight_rom[4837] = -42;
        weight_rom[4838] = -43;
        weight_rom[4839] = -55;
        weight_rom[4840] = -58;
        weight_rom[4841] = -3;
        weight_rom[4842] = 16;
        weight_rom[4843] = 3;
        weight_rom[4844] = 2;
        weight_rom[4845] = -2;
        weight_rom[4846] = 0;
        weight_rom[4847] = 23;
        weight_rom[4848] = 15;
        weight_rom[4849] = -1;
        weight_rom[4850] = 4;
        weight_rom[4851] = -4;
        weight_rom[4852] = 4;
        weight_rom[4853] = -3;
        weight_rom[4854] = -3;
        weight_rom[4855] = 15;
        weight_rom[4856] = 21;
        weight_rom[4857] = 32;
        weight_rom[4858] = 16;
        weight_rom[4859] = 22;
        weight_rom[4860] = 17;
        weight_rom[4861] = 15;
        weight_rom[4862] = 10;
        weight_rom[4863] = -2;
        weight_rom[4864] = -10;
        weight_rom[4865] = -10;
        weight_rom[4866] = -14;
        weight_rom[4867] = -42;
        weight_rom[4868] = -53;
        weight_rom[4869] = -25;
        weight_rom[4870] = -20;
        weight_rom[4871] = -4;
        weight_rom[4872] = 0;
        weight_rom[4873] = 2;
        weight_rom[4874] = 8;
        weight_rom[4875] = 38;
        weight_rom[4876] = 2;
        weight_rom[4877] = -12;
        weight_rom[4878] = 6;
        weight_rom[4879] = -10;
        weight_rom[4880] = -4;
        weight_rom[4881] = 9;
        weight_rom[4882] = 23;
        weight_rom[4883] = 27;
        weight_rom[4884] = 25;
        weight_rom[4885] = 45;
        weight_rom[4886] = 51;
        weight_rom[4887] = 37;
        weight_rom[4888] = 44;
        weight_rom[4889] = 34;
        weight_rom[4890] = 53;
        weight_rom[4891] = 22;
        weight_rom[4892] = 13;
        weight_rom[4893] = 7;
        weight_rom[4894] = -7;
        weight_rom[4895] = -41;
        weight_rom[4896] = -54;
        weight_rom[4897] = -48;
        weight_rom[4898] = -46;
        weight_rom[4899] = -15;
        weight_rom[4900] = -2;
        weight_rom[4901] = 16;
        weight_rom[4902] = 18;
        weight_rom[4903] = 38;
        weight_rom[4904] = 9;
        weight_rom[4905] = -5;
        weight_rom[4906] = 5;
        weight_rom[4907] = -6;
        weight_rom[4908] = 3;
        weight_rom[4909] = 14;
        weight_rom[4910] = 14;
        weight_rom[4911] = 19;
        weight_rom[4912] = 39;
        weight_rom[4913] = 42;
        weight_rom[4914] = 52;
        weight_rom[4915] = 48;
        weight_rom[4916] = 47;
        weight_rom[4917] = 46;
        weight_rom[4918] = 42;
        weight_rom[4919] = 37;
        weight_rom[4920] = 23;
        weight_rom[4921] = 14;
        weight_rom[4922] = 5;
        weight_rom[4923] = -13;
        weight_rom[4924] = -44;
        weight_rom[4925] = -60;
        weight_rom[4926] = -33;
        weight_rom[4927] = 7;
        weight_rom[4928] = 7;
        weight_rom[4929] = 11;
        weight_rom[4930] = 3;
        weight_rom[4931] = 16;
        weight_rom[4932] = 6;
        weight_rom[4933] = -9;
        weight_rom[4934] = 0;
        weight_rom[4935] = -3;
        weight_rom[4936] = 7;
        weight_rom[4937] = -1;
        weight_rom[4938] = 13;
        weight_rom[4939] = 11;
        weight_rom[4940] = 18;
        weight_rom[4941] = 33;
        weight_rom[4942] = 59;
        weight_rom[4943] = 55;
        weight_rom[4944] = 58;
        weight_rom[4945] = 53;
        weight_rom[4946] = 53;
        weight_rom[4947] = 43;
        weight_rom[4948] = 29;
        weight_rom[4949] = 20;
        weight_rom[4950] = 20;
        weight_rom[4951] = -7;
        weight_rom[4952] = -43;
        weight_rom[4953] = -51;
        weight_rom[4954] = -13;
        weight_rom[4955] = -16;
        weight_rom[4956] = 14;
        weight_rom[4957] = 13;
        weight_rom[4958] = 1;
        weight_rom[4959] = 20;
        weight_rom[4960] = 7;
        weight_rom[4961] = -6;
        weight_rom[4962] = -1;
        weight_rom[4963] = -6;
        weight_rom[4964] = -11;
        weight_rom[4965] = -6;
        weight_rom[4966] = -1;
        weight_rom[4967] = -10;
        weight_rom[4968] = 5;
        weight_rom[4969] = 25;
        weight_rom[4970] = 52;
        weight_rom[4971] = 56;
        weight_rom[4972] = 49;
        weight_rom[4973] = 56;
        weight_rom[4974] = 54;
        weight_rom[4975] = 40;
        weight_rom[4976] = 27;
        weight_rom[4977] = 9;
        weight_rom[4978] = 23;
        weight_rom[4979] = -10;
        weight_rom[4980] = -39;
        weight_rom[4981] = -37;
        weight_rom[4982] = -12;
        weight_rom[4983] = 11;
        weight_rom[4984] = 9;
        weight_rom[4985] = 14;
        weight_rom[4986] = 10;
        weight_rom[4987] = 28;
        weight_rom[4988] = -16;
        weight_rom[4989] = 1;
        weight_rom[4990] = 7;
        weight_rom[4991] = -15;
        weight_rom[4992] = -21;
        weight_rom[4993] = -27;
        weight_rom[4994] = -26;
        weight_rom[4995] = -29;
        weight_rom[4996] = -30;
        weight_rom[4997] = -9;
        weight_rom[4998] = 35;
        weight_rom[4999] = 28;
        weight_rom[5000] = 42;
        weight_rom[5001] = 47;
        weight_rom[5002] = 45;
        weight_rom[5003] = 34;
        weight_rom[5004] = 33;
        weight_rom[5005] = 21;
        weight_rom[5006] = 31;
        weight_rom[5007] = 18;
        weight_rom[5008] = -16;
        weight_rom[5009] = -44;
        weight_rom[5010] = -17;
        weight_rom[5011] = 1;
        weight_rom[5012] = 11;
        weight_rom[5013] = 14;
        weight_rom[5014] = 20;
        weight_rom[5015] = 16;
        weight_rom[5016] = -14;
        weight_rom[5017] = -24;
        weight_rom[5018] = -20;
        weight_rom[5019] = -19;
        weight_rom[5020] = -21;
        weight_rom[5021] = -40;
        weight_rom[5022] = -42;
        weight_rom[5023] = -38;
        weight_rom[5024] = -54;
        weight_rom[5025] = -30;
        weight_rom[5026] = -2;
        weight_rom[5027] = -3;
        weight_rom[5028] = -8;
        weight_rom[5029] = 17;
        weight_rom[5030] = 32;
        weight_rom[5031] = 25;
        weight_rom[5032] = 38;
        weight_rom[5033] = 38;
        weight_rom[5034] = 48;
        weight_rom[5035] = 11;
        weight_rom[5036] = -23;
        weight_rom[5037] = -8;
        weight_rom[5038] = -27;
        weight_rom[5039] = -5;
        weight_rom[5040] = 11;
        weight_rom[5041] = 1;
        weight_rom[5042] = 9;
        weight_rom[5043] = 3;
        weight_rom[5044] = -25;
        weight_rom[5045] = -20;
        weight_rom[5046] = -34;
        weight_rom[5047] = -37;
        weight_rom[5048] = -38;
        weight_rom[5049] = -34;
        weight_rom[5050] = -34;
        weight_rom[5051] = -47;
        weight_rom[5052] = -51;
        weight_rom[5053] = -40;
        weight_rom[5054] = -8;
        weight_rom[5055] = -9;
        weight_rom[5056] = -10;
        weight_rom[5057] = 1;
        weight_rom[5058] = 16;
        weight_rom[5059] = 27;
        weight_rom[5060] = 28;
        weight_rom[5061] = 14;
        weight_rom[5062] = 19;
        weight_rom[5063] = 2;
        weight_rom[5064] = 3;
        weight_rom[5065] = 7;
        weight_rom[5066] = -4;
        weight_rom[5067] = -8;
        weight_rom[5068] = -2;
        weight_rom[5069] = -4;
        weight_rom[5070] = 19;
        weight_rom[5071] = 5;
        weight_rom[5072] = -26;
        weight_rom[5073] = -36;
        weight_rom[5074] = -33;
        weight_rom[5075] = -33;
        weight_rom[5076] = -20;
        weight_rom[5077] = -21;
        weight_rom[5078] = -25;
        weight_rom[5079] = -30;
        weight_rom[5080] = -38;
        weight_rom[5081] = -18;
        weight_rom[5082] = -7;
        weight_rom[5083] = -17;
        weight_rom[5084] = -3;
        weight_rom[5085] = 3;
        weight_rom[5086] = 4;
        weight_rom[5087] = 10;
        weight_rom[5088] = -3;
        weight_rom[5089] = 1;
        weight_rom[5090] = -3;
        weight_rom[5091] = -6;
        weight_rom[5092] = 11;
        weight_rom[5093] = 7;
        weight_rom[5094] = 4;
        weight_rom[5095] = 14;
        weight_rom[5096] = -2;
        weight_rom[5097] = 5;
        weight_rom[5098] = 0;
        weight_rom[5099] = -1;
        weight_rom[5100] = -28;
        weight_rom[5101] = -28;
        weight_rom[5102] = -17;
        weight_rom[5103] = -7;
        weight_rom[5104] = -15;
        weight_rom[5105] = -15;
        weight_rom[5106] = -17;
        weight_rom[5107] = -27;
        weight_rom[5108] = -19;
        weight_rom[5109] = -5;
        weight_rom[5110] = -11;
        weight_rom[5111] = -9;
        weight_rom[5112] = -16;
        weight_rom[5113] = -6;
        weight_rom[5114] = 7;
        weight_rom[5115] = 6;
        weight_rom[5116] = 0;
        weight_rom[5117] = 0;
        weight_rom[5118] = -12;
        weight_rom[5119] = 0;
        weight_rom[5120] = 6;
        weight_rom[5121] = 4;
        weight_rom[5122] = 22;
        weight_rom[5123] = -4;
        weight_rom[5124] = -4;
        weight_rom[5125] = 3;
        weight_rom[5126] = 5;
        weight_rom[5127] = -3;
        weight_rom[5128] = 16;
        weight_rom[5129] = 7;
        weight_rom[5130] = -4;
        weight_rom[5131] = 3;
        weight_rom[5132] = -11;
        weight_rom[5133] = -13;
        weight_rom[5134] = -9;
        weight_rom[5135] = -14;
        weight_rom[5136] = -19;
        weight_rom[5137] = -15;
        weight_rom[5138] = -18;
        weight_rom[5139] = -14;
        weight_rom[5140] = -19;
        weight_rom[5141] = -4;
        weight_rom[5142] = 1;
        weight_rom[5143] = -3;
        weight_rom[5144] = -5;
        weight_rom[5145] = -6;
        weight_rom[5146] = -11;
        weight_rom[5147] = -6;
        weight_rom[5148] = 25;
        weight_rom[5149] = 8;
        weight_rom[5150] = 19;
        weight_rom[5151] = 14;
        weight_rom[5152] = -2;
        weight_rom[5153] = 2;
        weight_rom[5154] = 21;
        weight_rom[5155] = 24;
        weight_rom[5156] = 36;
        weight_rom[5157] = 22;
        weight_rom[5158] = 2;
        weight_rom[5159] = -6;
        weight_rom[5160] = -19;
        weight_rom[5161] = -2;
        weight_rom[5162] = -2;
        weight_rom[5163] = -9;
        weight_rom[5164] = -10;
        weight_rom[5165] = -15;
        weight_rom[5166] = -27;
        weight_rom[5167] = -25;
        weight_rom[5168] = -11;
        weight_rom[5169] = 2;
        weight_rom[5170] = -7;
        weight_rom[5171] = -7;
        weight_rom[5172] = -15;
        weight_rom[5173] = -2;
        weight_rom[5174] = -2;
        weight_rom[5175] = -1;
        weight_rom[5176] = 13;
        weight_rom[5177] = 19;
        weight_rom[5178] = 20;
        weight_rom[5179] = 22;
        weight_rom[5180] = 3;
        weight_rom[5181] = 15;
        weight_rom[5182] = 1;
        weight_rom[5183] = 40;
        weight_rom[5184] = 43;
        weight_rom[5185] = 13;
        weight_rom[5186] = 3;
        weight_rom[5187] = -5;
        weight_rom[5188] = -13;
        weight_rom[5189] = -10;
        weight_rom[5190] = -4;
        weight_rom[5191] = -6;
        weight_rom[5192] = -7;
        weight_rom[5193] = -21;
        weight_rom[5194] = -23;
        weight_rom[5195] = -11;
        weight_rom[5196] = -15;
        weight_rom[5197] = -4;
        weight_rom[5198] = -3;
        weight_rom[5199] = -4;
        weight_rom[5200] = -19;
        weight_rom[5201] = -18;
        weight_rom[5202] = -6;
        weight_rom[5203] = 7;
        weight_rom[5204] = 17;
        weight_rom[5205] = 40;
        weight_rom[5206] = 37;
        weight_rom[5207] = -2;
        weight_rom[5208] = -4;
        weight_rom[5209] = 13;
        weight_rom[5210] = 23;
        weight_rom[5211] = 18;
        weight_rom[5212] = 30;
        weight_rom[5213] = 22;
        weight_rom[5214] = 7;
        weight_rom[5215] = 1;
        weight_rom[5216] = -3;
        weight_rom[5217] = 0;
        weight_rom[5218] = 2;
        weight_rom[5219] = 1;
        weight_rom[5220] = -16;
        weight_rom[5221] = -14;
        weight_rom[5222] = -16;
        weight_rom[5223] = 0;
        weight_rom[5224] = 3;
        weight_rom[5225] = 12;
        weight_rom[5226] = 9;
        weight_rom[5227] = 4;
        weight_rom[5228] = -16;
        weight_rom[5229] = -14;
        weight_rom[5230] = 5;
        weight_rom[5231] = 11;
        weight_rom[5232] = 24;
        weight_rom[5233] = 44;
        weight_rom[5234] = 14;
        weight_rom[5235] = 17;
        weight_rom[5236] = -2;
        weight_rom[5237] = 16;
        weight_rom[5238] = -9;
        weight_rom[5239] = 17;
        weight_rom[5240] = 25;
        weight_rom[5241] = 17;
        weight_rom[5242] = 10;
        weight_rom[5243] = 14;
        weight_rom[5244] = 20;
        weight_rom[5245] = 15;
        weight_rom[5246] = 11;
        weight_rom[5247] = 1;
        weight_rom[5248] = 4;
        weight_rom[5249] = 7;
        weight_rom[5250] = 8;
        weight_rom[5251] = 0;
        weight_rom[5252] = 5;
        weight_rom[5253] = 15;
        weight_rom[5254] = -5;
        weight_rom[5255] = 2;
        weight_rom[5256] = -1;
        weight_rom[5257] = 1;
        weight_rom[5258] = 7;
        weight_rom[5259] = 14;
        weight_rom[5260] = 5;
        weight_rom[5261] = 31;
        weight_rom[5262] = 20;
        weight_rom[5263] = 9;
        weight_rom[5264] = 3;
        weight_rom[5265] = 15;
        weight_rom[5266] = -6;
        weight_rom[5267] = 18;
        weight_rom[5268] = 32;
        weight_rom[5269] = 36;
        weight_rom[5270] = 29;
        weight_rom[5271] = 23;
        weight_rom[5272] = 26;
        weight_rom[5273] = 13;
        weight_rom[5274] = 18;
        weight_rom[5275] = 10;
        weight_rom[5276] = 11;
        weight_rom[5277] = 9;
        weight_rom[5278] = 10;
        weight_rom[5279] = 5;
        weight_rom[5280] = 6;
        weight_rom[5281] = -2;
        weight_rom[5282] = -10;
        weight_rom[5283] = -6;
        weight_rom[5284] = -10;
        weight_rom[5285] = 0;
        weight_rom[5286] = -3;
        weight_rom[5287] = 1;
        weight_rom[5288] = 14;
        weight_rom[5289] = 7;
        weight_rom[5290] = 7;
        weight_rom[5291] = -1;
        weight_rom[5292] = 2;
        weight_rom[5293] = 19;
        weight_rom[5294] = 40;
        weight_rom[5295] = 39;
        weight_rom[5296] = 27;
        weight_rom[5297] = 24;
        weight_rom[5298] = 36;
        weight_rom[5299] = 31;
        weight_rom[5300] = 21;
        weight_rom[5301] = 19;
        weight_rom[5302] = 18;
        weight_rom[5303] = 19;
        weight_rom[5304] = 6;
        weight_rom[5305] = 1;
        weight_rom[5306] = 7;
        weight_rom[5307] = 0;
        weight_rom[5308] = 5;
        weight_rom[5309] = -12;
        weight_rom[5310] = 4;
        weight_rom[5311] = -1;
        weight_rom[5312] = -14;
        weight_rom[5313] = 5;
        weight_rom[5314] = -9;
        weight_rom[5315] = 8;
        weight_rom[5316] = 21;
        weight_rom[5317] = 19;
        weight_rom[5318] = -5;
        weight_rom[5319] = 3;
        weight_rom[5320] = 4;
        weight_rom[5321] = -1;
        weight_rom[5322] = 32;
        weight_rom[5323] = 39;
        weight_rom[5324] = 13;
        weight_rom[5325] = 26;
        weight_rom[5326] = 47;
        weight_rom[5327] = 34;
        weight_rom[5328] = 37;
        weight_rom[5329] = 38;
        weight_rom[5330] = 22;
        weight_rom[5331] = 24;
        weight_rom[5332] = 13;
        weight_rom[5333] = 8;
        weight_rom[5334] = 12;
        weight_rom[5335] = 8;
        weight_rom[5336] = 8;
        weight_rom[5337] = -2;
        weight_rom[5338] = -11;
        weight_rom[5339] = -3;
        weight_rom[5340] = -10;
        weight_rom[5341] = -20;
        weight_rom[5342] = 16;
        weight_rom[5343] = 9;
        weight_rom[5344] = 21;
        weight_rom[5345] = 9;
        weight_rom[5346] = 1;
        weight_rom[5347] = 2;
        weight_rom[5348] = -2;
        weight_rom[5349] = 2;
        weight_rom[5350] = 16;
        weight_rom[5351] = 18;
        weight_rom[5352] = 15;
        weight_rom[5353] = 23;
        weight_rom[5354] = 35;
        weight_rom[5355] = 49;
        weight_rom[5356] = 38;
        weight_rom[5357] = 29;
        weight_rom[5358] = 32;
        weight_rom[5359] = 30;
        weight_rom[5360] = 20;
        weight_rom[5361] = 15;
        weight_rom[5362] = 9;
        weight_rom[5363] = 5;
        weight_rom[5364] = -7;
        weight_rom[5365] = -2;
        weight_rom[5366] = -5;
        weight_rom[5367] = -21;
        weight_rom[5368] = -26;
        weight_rom[5369] = -9;
        weight_rom[5370] = 21;
        weight_rom[5371] = 16;
        weight_rom[5372] = 21;
        weight_rom[5373] = -9;
        weight_rom[5374] = 12;
        weight_rom[5375] = 4;
        weight_rom[5376] = 3;
        weight_rom[5377] = -1;
        weight_rom[5378] = 2;
        weight_rom[5379] = 16;
        weight_rom[5380] = 49;
        weight_rom[5381] = 54;
        weight_rom[5382] = 32;
        weight_rom[5383] = 24;
        weight_rom[5384] = 12;
        weight_rom[5385] = 4;
        weight_rom[5386] = 14;
        weight_rom[5387] = 7;
        weight_rom[5388] = 15;
        weight_rom[5389] = 19;
        weight_rom[5390] = 10;
        weight_rom[5391] = 8;
        weight_rom[5392] = 5;
        weight_rom[5393] = 24;
        weight_rom[5394] = -5;
        weight_rom[5395] = -14;
        weight_rom[5396] = -7;
        weight_rom[5397] = 22;
        weight_rom[5398] = 17;
        weight_rom[5399] = 11;
        weight_rom[5400] = 20;
        weight_rom[5401] = 24;
        weight_rom[5402] = 3;
        weight_rom[5403] = 3;
        weight_rom[5404] = 1;
        weight_rom[5405] = 4;
        weight_rom[5406] = -2;
        weight_rom[5407] = -10;
        weight_rom[5408] = 12;
        weight_rom[5409] = 38;
        weight_rom[5410] = 25;
        weight_rom[5411] = 36;
        weight_rom[5412] = 53;
        weight_rom[5413] = 38;
        weight_rom[5414] = 14;
        weight_rom[5415] = 30;
        weight_rom[5416] = 35;
        weight_rom[5417] = 31;
        weight_rom[5418] = 22;
        weight_rom[5419] = 23;
        weight_rom[5420] = 26;
        weight_rom[5421] = 22;
        weight_rom[5422] = 31;
        weight_rom[5423] = 27;
        weight_rom[5424] = 22;
        weight_rom[5425] = 48;
        weight_rom[5426] = 10;
        weight_rom[5427] = 1;
        weight_rom[5428] = 0;
        weight_rom[5429] = -2;
        weight_rom[5430] = -3;
        weight_rom[5431] = 1;
        weight_rom[5432] = -4;
        weight_rom[5433] = -2;
        weight_rom[5434] = -1;
        weight_rom[5435] = 2;
        weight_rom[5436] = 23;
        weight_rom[5437] = 7;
        weight_rom[5438] = 20;
        weight_rom[5439] = 58;
        weight_rom[5440] = 60;
        weight_rom[5441] = 60;
        weight_rom[5442] = 53;
        weight_rom[5443] = 46;
        weight_rom[5444] = 31;
        weight_rom[5445] = 65;
        weight_rom[5446] = 76;
        weight_rom[5447] = 48;
        weight_rom[5448] = 66;
        weight_rom[5449] = 65;
        weight_rom[5450] = 60;
        weight_rom[5451] = 53;
        weight_rom[5452] = 40;
        weight_rom[5453] = 30;
        weight_rom[5454] = 34;
        weight_rom[5455] = 17;
        weight_rom[5456] = 0;
        weight_rom[5457] = 3;
        weight_rom[5458] = -3;
        weight_rom[5459] = -3;
        weight_rom[5460] = -3;
        weight_rom[5461] = 4;
        weight_rom[5462] = 0;
        weight_rom[5463] = 4;
        weight_rom[5464] = 1;
        weight_rom[5465] = 13;
        weight_rom[5466] = 6;
        weight_rom[5467] = 19;
        weight_rom[5468] = 27;
        weight_rom[5469] = 22;
        weight_rom[5470] = 33;
        weight_rom[5471] = 16;
        weight_rom[5472] = 23;
        weight_rom[5473] = 24;
        weight_rom[5474] = 43;
        weight_rom[5475] = 32;
        weight_rom[5476] = 28;
        weight_rom[5477] = 33;
        weight_rom[5478] = 40;
        weight_rom[5479] = 24;
        weight_rom[5480] = 18;
        weight_rom[5481] = 2;
        weight_rom[5482] = 11;
        weight_rom[5483] = 4;
        weight_rom[5484] = 2;
        weight_rom[5485] = -2;
        weight_rom[5486] = -2;
        weight_rom[5487] = 0;
        weight_rom[5488] = -2;
        weight_rom[5489] = 0;
        weight_rom[5490] = 1;
        weight_rom[5491] = -1;
        weight_rom[5492] = 1;
        weight_rom[5493] = 0;
        weight_rom[5494] = 2;
        weight_rom[5495] = -1;
        weight_rom[5496] = -2;
        weight_rom[5497] = -1;
        weight_rom[5498] = -3;
        weight_rom[5499] = -3;
        weight_rom[5500] = -4;
        weight_rom[5501] = -9;
        weight_rom[5502] = 3;
        weight_rom[5503] = -4;
        weight_rom[5504] = 4;
        weight_rom[5505] = 4;
        weight_rom[5506] = 2;
        weight_rom[5507] = -2;
        weight_rom[5508] = -3;
        weight_rom[5509] = -4;
        weight_rom[5510] = 3;
        weight_rom[5511] = -1;
        weight_rom[5512] = 4;
        weight_rom[5513] = 0;
        weight_rom[5514] = 3;
        weight_rom[5515] = -2;
        weight_rom[5516] = -3;
        weight_rom[5517] = -4;
        weight_rom[5518] = 1;
        weight_rom[5519] = 0;
        weight_rom[5520] = 3;
        weight_rom[5521] = -4;
        weight_rom[5522] = -6;
        weight_rom[5523] = -3;
        weight_rom[5524] = -7;
        weight_rom[5525] = -6;
        weight_rom[5526] = 1;
        weight_rom[5527] = 0;
        weight_rom[5528] = -9;
        weight_rom[5529] = -19;
        weight_rom[5530] = 8;
        weight_rom[5531] = 9;
        weight_rom[5532] = 2;
        weight_rom[5533] = -8;
        weight_rom[5534] = -6;
        weight_rom[5535] = -7;
        weight_rom[5536] = 0;
        weight_rom[5537] = 4;
        weight_rom[5538] = -4;
        weight_rom[5539] = 1;
        weight_rom[5540] = 1;
        weight_rom[5541] = -1;
        weight_rom[5542] = -2;
        weight_rom[5543] = -2;
        weight_rom[5544] = -4;
        weight_rom[5545] = 1;
        weight_rom[5546] = 2;
        weight_rom[5547] = 2;
        weight_rom[5548] = -2;
        weight_rom[5549] = -3;
        weight_rom[5550] = -7;
        weight_rom[5551] = -17;
        weight_rom[5552] = -11;
        weight_rom[5553] = -6;
        weight_rom[5554] = -29;
        weight_rom[5555] = -23;
        weight_rom[5556] = -43;
        weight_rom[5557] = -31;
        weight_rom[5558] = -40;
        weight_rom[5559] = -4;
        weight_rom[5560] = 2;
        weight_rom[5561] = -3;
        weight_rom[5562] = -4;
        weight_rom[5563] = 14;
        weight_rom[5564] = -8;
        weight_rom[5565] = 3;
        weight_rom[5566] = 3;
        weight_rom[5567] = -9;
        weight_rom[5568] = -2;
        weight_rom[5569] = 3;
        weight_rom[5570] = 1;
        weight_rom[5571] = 1;
        weight_rom[5572] = 1;
        weight_rom[5573] = -4;
        weight_rom[5574] = -1;
        weight_rom[5575] = 3;
        weight_rom[5576] = 4;
        weight_rom[5577] = 19;
        weight_rom[5578] = 17;
        weight_rom[5579] = 22;
        weight_rom[5580] = 25;
        weight_rom[5581] = 5;
        weight_rom[5582] = 14;
        weight_rom[5583] = 16;
        weight_rom[5584] = 10;
        weight_rom[5585] = 0;
        weight_rom[5586] = 17;
        weight_rom[5587] = 8;
        weight_rom[5588] = 3;
        weight_rom[5589] = 17;
        weight_rom[5590] = 9;
        weight_rom[5591] = 14;
        weight_rom[5592] = 28;
        weight_rom[5593] = 1;
        weight_rom[5594] = 7;
        weight_rom[5595] = 2;
        weight_rom[5596] = -7;
        weight_rom[5597] = -4;
        weight_rom[5598] = -4;
        weight_rom[5599] = 3;
        weight_rom[5600] = 1;
        weight_rom[5601] = -4;
        weight_rom[5602] = 14;
        weight_rom[5603] = 3;
        weight_rom[5604] = 15;
        weight_rom[5605] = 27;
        weight_rom[5606] = 28;
        weight_rom[5607] = 24;
        weight_rom[5608] = 29;
        weight_rom[5609] = 15;
        weight_rom[5610] = 18;
        weight_rom[5611] = 31;
        weight_rom[5612] = 26;
        weight_rom[5613] = 16;
        weight_rom[5614] = 9;
        weight_rom[5615] = 10;
        weight_rom[5616] = 17;
        weight_rom[5617] = 2;
        weight_rom[5618] = 16;
        weight_rom[5619] = 5;
        weight_rom[5620] = -5;
        weight_rom[5621] = 5;
        weight_rom[5622] = 2;
        weight_rom[5623] = -11;
        weight_rom[5624] = 16;
        weight_rom[5625] = 7;
        weight_rom[5626] = 12;
        weight_rom[5627] = 1;
        weight_rom[5628] = -4;
        weight_rom[5629] = 3;
        weight_rom[5630] = -1;
        weight_rom[5631] = 5;
        weight_rom[5632] = 13;
        weight_rom[5633] = 27;
        weight_rom[5634] = 15;
        weight_rom[5635] = 15;
        weight_rom[5636] = -5;
        weight_rom[5637] = 9;
        weight_rom[5638] = 13;
        weight_rom[5639] = 24;
        weight_rom[5640] = 25;
        weight_rom[5641] = 16;
        weight_rom[5642] = 8;
        weight_rom[5643] = 3;
        weight_rom[5644] = 3;
        weight_rom[5645] = -5;
        weight_rom[5646] = -7;
        weight_rom[5647] = -9;
        weight_rom[5648] = 0;
        weight_rom[5649] = -11;
        weight_rom[5650] = 5;
        weight_rom[5651] = -3;
        weight_rom[5652] = -5;
        weight_rom[5653] = 21;
        weight_rom[5654] = 3;
        weight_rom[5655] = 0;
        weight_rom[5656] = 0;
        weight_rom[5657] = -1;
        weight_rom[5658] = 7;
        weight_rom[5659] = 2;
        weight_rom[5660] = 20;
        weight_rom[5661] = 6;
        weight_rom[5662] = -7;
        weight_rom[5663] = -3;
        weight_rom[5664] = -1;
        weight_rom[5665] = 3;
        weight_rom[5666] = 10;
        weight_rom[5667] = 17;
        weight_rom[5668] = 9;
        weight_rom[5669] = 20;
        weight_rom[5670] = 12;
        weight_rom[5671] = 10;
        weight_rom[5672] = 17;
        weight_rom[5673] = 5;
        weight_rom[5674] = 11;
        weight_rom[5675] = 0;
        weight_rom[5676] = 5;
        weight_rom[5677] = -3;
        weight_rom[5678] = -1;
        weight_rom[5679] = -4;
        weight_rom[5680] = 8;
        weight_rom[5681] = 5;
        weight_rom[5682] = 3;
        weight_rom[5683] = 0;
        weight_rom[5684] = -4;
        weight_rom[5685] = 8;
        weight_rom[5686] = -22;
        weight_rom[5687] = -1;
        weight_rom[5688] = -8;
        weight_rom[5689] = 8;
        weight_rom[5690] = -2;
        weight_rom[5691] = -19;
        weight_rom[5692] = -5;
        weight_rom[5693] = -6;
        weight_rom[5694] = -4;
        weight_rom[5695] = 3;
        weight_rom[5696] = 10;
        weight_rom[5697] = 11;
        weight_rom[5698] = 23;
        weight_rom[5699] = 23;
        weight_rom[5700] = 12;
        weight_rom[5701] = 7;
        weight_rom[5702] = 0;
        weight_rom[5703] = 2;
        weight_rom[5704] = 1;
        weight_rom[5705] = 4;
        weight_rom[5706] = -23;
        weight_rom[5707] = -25;
        weight_rom[5708] = -3;
        weight_rom[5709] = 16;
        weight_rom[5710] = -7;
        weight_rom[5711] = -4;
        weight_rom[5712] = -3;
        weight_rom[5713] = -6;
        weight_rom[5714] = -6;
        weight_rom[5715] = -22;
        weight_rom[5716] = -12;
        weight_rom[5717] = -1;
        weight_rom[5718] = -15;
        weight_rom[5719] = -13;
        weight_rom[5720] = -3;
        weight_rom[5721] = 1;
        weight_rom[5722] = -3;
        weight_rom[5723] = 4;
        weight_rom[5724] = -15;
        weight_rom[5725] = 4;
        weight_rom[5726] = 16;
        weight_rom[5727] = 7;
        weight_rom[5728] = -3;
        weight_rom[5729] = -13;
        weight_rom[5730] = -23;
        weight_rom[5731] = -10;
        weight_rom[5732] = -12;
        weight_rom[5733] = -1;
        weight_rom[5734] = -20;
        weight_rom[5735] = -33;
        weight_rom[5736] = -12;
        weight_rom[5737] = 28;
        weight_rom[5738] = 4;
        weight_rom[5739] = -6;
        weight_rom[5740] = -1;
        weight_rom[5741] = -4;
        weight_rom[5742] = -9;
        weight_rom[5743] = -14;
        weight_rom[5744] = -13;
        weight_rom[5745] = -11;
        weight_rom[5746] = -8;
        weight_rom[5747] = 3;
        weight_rom[5748] = 0;
        weight_rom[5749] = 5;
        weight_rom[5750] = -1;
        weight_rom[5751] = 0;
        weight_rom[5752] = -4;
        weight_rom[5753] = 2;
        weight_rom[5754] = 0;
        weight_rom[5755] = 8;
        weight_rom[5756] = -24;
        weight_rom[5757] = -38;
        weight_rom[5758] = -28;
        weight_rom[5759] = -27;
        weight_rom[5760] = -20;
        weight_rom[5761] = -10;
        weight_rom[5762] = 10;
        weight_rom[5763] = -24;
        weight_rom[5764] = 0;
        weight_rom[5765] = 21;
        weight_rom[5766] = 3;
        weight_rom[5767] = 1;
        weight_rom[5768] = -5;
        weight_rom[5769] = -9;
        weight_rom[5770] = -27;
        weight_rom[5771] = -11;
        weight_rom[5772] = -24;
        weight_rom[5773] = -28;
        weight_rom[5774] = -11;
        weight_rom[5775] = 2;
        weight_rom[5776] = 21;
        weight_rom[5777] = -1;
        weight_rom[5778] = 5;
        weight_rom[5779] = 10;
        weight_rom[5780] = 5;
        weight_rom[5781] = -3;
        weight_rom[5782] = -6;
        weight_rom[5783] = -11;
        weight_rom[5784] = -29;
        weight_rom[5785] = -27;
        weight_rom[5786] = -28;
        weight_rom[5787] = -31;
        weight_rom[5788] = -25;
        weight_rom[5789] = -25;
        weight_rom[5790] = -22;
        weight_rom[5791] = -16;
        weight_rom[5792] = -1;
        weight_rom[5793] = 35;
        weight_rom[5794] = 23;
        weight_rom[5795] = -1;
        weight_rom[5796] = 2;
        weight_rom[5797] = -15;
        weight_rom[5798] = -38;
        weight_rom[5799] = -18;
        weight_rom[5800] = -23;
        weight_rom[5801] = -9;
        weight_rom[5802] = -10;
        weight_rom[5803] = -7;
        weight_rom[5804] = 10;
        weight_rom[5805] = 7;
        weight_rom[5806] = 8;
        weight_rom[5807] = 22;
        weight_rom[5808] = 20;
        weight_rom[5809] = 23;
        weight_rom[5810] = 25;
        weight_rom[5811] = 12;
        weight_rom[5812] = 1;
        weight_rom[5813] = 9;
        weight_rom[5814] = 0;
        weight_rom[5815] = -2;
        weight_rom[5816] = -15;
        weight_rom[5817] = -24;
        weight_rom[5818] = -37;
        weight_rom[5819] = -33;
        weight_rom[5820] = -18;
        weight_rom[5821] = 15;
        weight_rom[5822] = 14;
        weight_rom[5823] = -2;
        weight_rom[5824] = 2;
        weight_rom[5825] = -11;
        weight_rom[5826] = -34;
        weight_rom[5827] = -43;
        weight_rom[5828] = -36;
        weight_rom[5829] = -15;
        weight_rom[5830] = -6;
        weight_rom[5831] = 0;
        weight_rom[5832] = -6;
        weight_rom[5833] = 7;
        weight_rom[5834] = 29;
        weight_rom[5835] = 29;
        weight_rom[5836] = 32;
        weight_rom[5837] = 41;
        weight_rom[5838] = 47;
        weight_rom[5839] = 30;
        weight_rom[5840] = 16;
        weight_rom[5841] = 18;
        weight_rom[5842] = 11;
        weight_rom[5843] = 9;
        weight_rom[5844] = 3;
        weight_rom[5845] = -21;
        weight_rom[5846] = -25;
        weight_rom[5847] = -34;
        weight_rom[5848] = -52;
        weight_rom[5849] = -15;
        weight_rom[5850] = 7;
        weight_rom[5851] = -3;
        weight_rom[5852] = -1;
        weight_rom[5853] = -8;
        weight_rom[5854] = -27;
        weight_rom[5855] = -49;
        weight_rom[5856] = -34;
        weight_rom[5857] = -12;
        weight_rom[5858] = -15;
        weight_rom[5859] = 4;
        weight_rom[5860] = 7;
        weight_rom[5861] = 17;
        weight_rom[5862] = 16;
        weight_rom[5863] = 28;
        weight_rom[5864] = 33;
        weight_rom[5865] = 45;
        weight_rom[5866] = 47;
        weight_rom[5867] = 33;
        weight_rom[5868] = 27;
        weight_rom[5869] = 14;
        weight_rom[5870] = 6;
        weight_rom[5871] = 0;
        weight_rom[5872] = -17;
        weight_rom[5873] = -8;
        weight_rom[5874] = -6;
        weight_rom[5875] = -27;
        weight_rom[5876] = -50;
        weight_rom[5877] = -35;
        weight_rom[5878] = -2;
        weight_rom[5879] = 3;
        weight_rom[5880] = 1;
        weight_rom[5881] = -6;
        weight_rom[5882] = -11;
        weight_rom[5883] = -38;
        weight_rom[5884] = -47;
        weight_rom[5885] = -33;
        weight_rom[5886] = -16;
        weight_rom[5887] = -13;
        weight_rom[5888] = 7;
        weight_rom[5889] = 12;
        weight_rom[5890] = 22;
        weight_rom[5891] = 17;
        weight_rom[5892] = 27;
        weight_rom[5893] = 28;
        weight_rom[5894] = 38;
        weight_rom[5895] = 24;
        weight_rom[5896] = 15;
        weight_rom[5897] = 3;
        weight_rom[5898] = -7;
        weight_rom[5899] = -23;
        weight_rom[5900] = -17;
        weight_rom[5901] = -8;
        weight_rom[5902] = -9;
        weight_rom[5903] = -5;
        weight_rom[5904] = -11;
        weight_rom[5905] = -11;
        weight_rom[5906] = -8;
        weight_rom[5907] = 2;
        weight_rom[5908] = -4;
        weight_rom[5909] = 7;
        weight_rom[5910] = 12;
        weight_rom[5911] = -24;
        weight_rom[5912] = -43;
        weight_rom[5913] = -54;
        weight_rom[5914] = -44;
        weight_rom[5915] = -46;
        weight_rom[5916] = -32;
        weight_rom[5917] = -2;
        weight_rom[5918] = 12;
        weight_rom[5919] = 35;
        weight_rom[5920] = 29;
        weight_rom[5921] = 23;
        weight_rom[5922] = 15;
        weight_rom[5923] = 7;
        weight_rom[5924] = 14;
        weight_rom[5925] = -12;
        weight_rom[5926] = -16;
        weight_rom[5927] = -10;
        weight_rom[5928] = -12;
        weight_rom[5929] = 0;
        weight_rom[5930] = 3;
        weight_rom[5931] = 14;
        weight_rom[5932] = 15;
        weight_rom[5933] = 2;
        weight_rom[5934] = 2;
        weight_rom[5935] = -9;
        weight_rom[5936] = -3;
        weight_rom[5937] = -3;
        weight_rom[5938] = 30;
        weight_rom[5939] = -10;
        weight_rom[5940] = -47;
        weight_rom[5941] = -65;
        weight_rom[5942] = -78;
        weight_rom[5943] = -90;
        weight_rom[5944] = -90;
        weight_rom[5945] = -58;
        weight_rom[5946] = -30;
        weight_rom[5947] = 12;
        weight_rom[5948] = 13;
        weight_rom[5949] = 9;
        weight_rom[5950] = -4;
        weight_rom[5951] = -14;
        weight_rom[5952] = -6;
        weight_rom[5953] = -25;
        weight_rom[5954] = -4;
        weight_rom[5955] = -6;
        weight_rom[5956] = -2;
        weight_rom[5957] = 3;
        weight_rom[5958] = 19;
        weight_rom[5959] = 22;
        weight_rom[5960] = 42;
        weight_rom[5961] = -14;
        weight_rom[5962] = -10;
        weight_rom[5963] = -1;
        weight_rom[5964] = -1;
        weight_rom[5965] = 7;
        weight_rom[5966] = 1;
        weight_rom[5967] = 13;
        weight_rom[5968] = -18;
        weight_rom[5969] = -32;
        weight_rom[5970] = -61;
        weight_rom[5971] = -80;
        weight_rom[5972] = -94;
        weight_rom[5973] = -127;
        weight_rom[5974] = -108;
        weight_rom[5975] = -93;
        weight_rom[5976] = -77;
        weight_rom[5977] = -61;
        weight_rom[5978] = -29;
        weight_rom[5979] = -6;
        weight_rom[5980] = -16;
        weight_rom[5981] = -9;
        weight_rom[5982] = -2;
        weight_rom[5983] = 4;
        weight_rom[5984] = 11;
        weight_rom[5985] = 29;
        weight_rom[5986] = 14;
        weight_rom[5987] = 23;
        weight_rom[5988] = 2;
        weight_rom[5989] = -33;
        weight_rom[5990] = -15;
        weight_rom[5991] = 2;
        weight_rom[5992] = -3;
        weight_rom[5993] = 8;
        weight_rom[5994] = 10;
        weight_rom[5995] = 41;
        weight_rom[5996] = 12;
        weight_rom[5997] = -18;
        weight_rom[5998] = -17;
        weight_rom[5999] = -52;
        weight_rom[6000] = -78;
        weight_rom[6001] = -101;
        weight_rom[6002] = -118;
        weight_rom[6003] = -122;
        weight_rom[6004] = -121;
        weight_rom[6005] = -68;
        weight_rom[6006] = -23;
        weight_rom[6007] = -8;
        weight_rom[6008] = -3;
        weight_rom[6009] = 2;
        weight_rom[6010] = 1;
        weight_rom[6011] = 20;
        weight_rom[6012] = 18;
        weight_rom[6013] = 28;
        weight_rom[6014] = 21;
        weight_rom[6015] = 21;
        weight_rom[6016] = 24;
        weight_rom[6017] = -3;
        weight_rom[6018] = -11;
        weight_rom[6019] = -5;
        weight_rom[6020] = 0;
        weight_rom[6021] = 6;
        weight_rom[6022] = 8;
        weight_rom[6023] = 57;
        weight_rom[6024] = 24;
        weight_rom[6025] = 17;
        weight_rom[6026] = 2;
        weight_rom[6027] = -10;
        weight_rom[6028] = -23;
        weight_rom[6029] = -31;
        weight_rom[6030] = -47;
        weight_rom[6031] = -54;
        weight_rom[6032] = -53;
        weight_rom[6033] = -26;
        weight_rom[6034] = -10;
        weight_rom[6035] = -5;
        weight_rom[6036] = 7;
        weight_rom[6037] = 4;
        weight_rom[6038] = 12;
        weight_rom[6039] = 10;
        weight_rom[6040] = 12;
        weight_rom[6041] = 25;
        weight_rom[6042] = 18;
        weight_rom[6043] = 22;
        weight_rom[6044] = 22;
        weight_rom[6045] = -6;
        weight_rom[6046] = -7;
        weight_rom[6047] = -8;
        weight_rom[6048] = 1;
        weight_rom[6049] = 7;
        weight_rom[6050] = 6;
        weight_rom[6051] = 45;
        weight_rom[6052] = 26;
        weight_rom[6053] = 18;
        weight_rom[6054] = 16;
        weight_rom[6055] = 14;
        weight_rom[6056] = 25;
        weight_rom[6057] = 26;
        weight_rom[6058] = 18;
        weight_rom[6059] = 6;
        weight_rom[6060] = -19;
        weight_rom[6061] = -7;
        weight_rom[6062] = 0;
        weight_rom[6063] = 4;
        weight_rom[6064] = 7;
        weight_rom[6065] = 14;
        weight_rom[6066] = 15;
        weight_rom[6067] = 13;
        weight_rom[6068] = 24;
        weight_rom[6069] = 13;
        weight_rom[6070] = 18;
        weight_rom[6071] = 22;
        weight_rom[6072] = 12;
        weight_rom[6073] = -15;
        weight_rom[6074] = -14;
        weight_rom[6075] = 3;
        weight_rom[6076] = 2;
        weight_rom[6077] = 5;
        weight_rom[6078] = 16;
        weight_rom[6079] = 24;
        weight_rom[6080] = 38;
        weight_rom[6081] = 24;
        weight_rom[6082] = 20;
        weight_rom[6083] = 18;
        weight_rom[6084] = 34;
        weight_rom[6085] = 31;
        weight_rom[6086] = 32;
        weight_rom[6087] = 8;
        weight_rom[6088] = 14;
        weight_rom[6089] = 3;
        weight_rom[6090] = 0;
        weight_rom[6091] = 2;
        weight_rom[6092] = 1;
        weight_rom[6093] = 5;
        weight_rom[6094] = 12;
        weight_rom[6095] = 15;
        weight_rom[6096] = 11;
        weight_rom[6097] = 14;
        weight_rom[6098] = 13;
        weight_rom[6099] = 15;
        weight_rom[6100] = -11;
        weight_rom[6101] = -26;
        weight_rom[6102] = -4;
        weight_rom[6103] = -3;
        weight_rom[6104] = -1;
        weight_rom[6105] = 4;
        weight_rom[6106] = 19;
        weight_rom[6107] = 34;
        weight_rom[6108] = 49;
        weight_rom[6109] = 15;
        weight_rom[6110] = -4;
        weight_rom[6111] = 7;
        weight_rom[6112] = 12;
        weight_rom[6113] = 22;
        weight_rom[6114] = 23;
        weight_rom[6115] = 15;
        weight_rom[6116] = 9;
        weight_rom[6117] = -2;
        weight_rom[6118] = 3;
        weight_rom[6119] = -1;
        weight_rom[6120] = 0;
        weight_rom[6121] = 7;
        weight_rom[6122] = 9;
        weight_rom[6123] = 3;
        weight_rom[6124] = 17;
        weight_rom[6125] = 1;
        weight_rom[6126] = -2;
        weight_rom[6127] = 5;
        weight_rom[6128] = -22;
        weight_rom[6129] = -23;
        weight_rom[6130] = 2;
        weight_rom[6131] = -4;
        weight_rom[6132] = 0;
        weight_rom[6133] = 3;
        weight_rom[6134] = 9;
        weight_rom[6135] = 51;
        weight_rom[6136] = 51;
        weight_rom[6137] = 32;
        weight_rom[6138] = 23;
        weight_rom[6139] = 16;
        weight_rom[6140] = 16;
        weight_rom[6141] = 12;
        weight_rom[6142] = 18;
        weight_rom[6143] = 5;
        weight_rom[6144] = 6;
        weight_rom[6145] = 4;
        weight_rom[6146] = -4;
        weight_rom[6147] = -5;
        weight_rom[6148] = -7;
        weight_rom[6149] = -1;
        weight_rom[6150] = -4;
        weight_rom[6151] = -12;
        weight_rom[6152] = -3;
        weight_rom[6153] = -7;
        weight_rom[6154] = -27;
        weight_rom[6155] = 0;
        weight_rom[6156] = 6;
        weight_rom[6157] = -12;
        weight_rom[6158] = 8;
        weight_rom[6159] = -1;
        weight_rom[6160] = 1;
        weight_rom[6161] = -3;
        weight_rom[6162] = 6;
        weight_rom[6163] = 21;
        weight_rom[6164] = 38;
        weight_rom[6165] = 36;
        weight_rom[6166] = 41;
        weight_rom[6167] = 43;
        weight_rom[6168] = 34;
        weight_rom[6169] = 30;
        weight_rom[6170] = 25;
        weight_rom[6171] = 23;
        weight_rom[6172] = 6;
        weight_rom[6173] = 5;
        weight_rom[6174] = -3;
        weight_rom[6175] = -3;
        weight_rom[6176] = -8;
        weight_rom[6177] = 1;
        weight_rom[6178] = -19;
        weight_rom[6179] = -33;
        weight_rom[6180] = -4;
        weight_rom[6181] = 4;
        weight_rom[6182] = 10;
        weight_rom[6183] = 18;
        weight_rom[6184] = 0;
        weight_rom[6185] = -2;
        weight_rom[6186] = 3;
        weight_rom[6187] = -2;
        weight_rom[6188] = -1;
        weight_rom[6189] = 4;
        weight_rom[6190] = 3;
        weight_rom[6191] = 6;
        weight_rom[6192] = 27;
        weight_rom[6193] = 32;
        weight_rom[6194] = 33;
        weight_rom[6195] = 44;
        weight_rom[6196] = 51;
        weight_rom[6197] = 47;
        weight_rom[6198] = 43;
        weight_rom[6199] = 28;
        weight_rom[6200] = 36;
        weight_rom[6201] = 19;
        weight_rom[6202] = 17;
        weight_rom[6203] = 7;
        weight_rom[6204] = 4;
        weight_rom[6205] = -6;
        weight_rom[6206] = -7;
        weight_rom[6207] = -4;
        weight_rom[6208] = 7;
        weight_rom[6209] = 14;
        weight_rom[6210] = 17;
        weight_rom[6211] = 26;
        weight_rom[6212] = 15;
        weight_rom[6213] = 1;
        weight_rom[6214] = 4;
        weight_rom[6215] = 2;
        weight_rom[6216] = -1;
        weight_rom[6217] = -2;
        weight_rom[6218] = 0;
        weight_rom[6219] = 3;
        weight_rom[6220] = 23;
        weight_rom[6221] = 20;
        weight_rom[6222] = 19;
        weight_rom[6223] = 27;
        weight_rom[6224] = 22;
        weight_rom[6225] = 31;
        weight_rom[6226] = 16;
        weight_rom[6227] = 16;
        weight_rom[6228] = 7;
        weight_rom[6229] = 14;
        weight_rom[6230] = 18;
        weight_rom[6231] = 10;
        weight_rom[6232] = 11;
        weight_rom[6233] = 3;
        weight_rom[6234] = 5;
        weight_rom[6235] = -15;
        weight_rom[6236] = -2;
        weight_rom[6237] = 2;
        weight_rom[6238] = 10;
        weight_rom[6239] = 4;
        weight_rom[6240] = -4;
        weight_rom[6241] = -1;
        weight_rom[6242] = 2;
        weight_rom[6243] = 0;
        weight_rom[6244] = 3;
        weight_rom[6245] = -3;
        weight_rom[6246] = 2;
        weight_rom[6247] = -2;
        weight_rom[6248] = 0;
        weight_rom[6249] = -6;
        weight_rom[6250] = -3;
        weight_rom[6251] = -6;
        weight_rom[6252] = -14;
        weight_rom[6253] = 8;
        weight_rom[6254] = -9;
        weight_rom[6255] = 8;
        weight_rom[6256] = 6;
        weight_rom[6257] = -22;
        weight_rom[6258] = 1;
        weight_rom[6259] = 19;
        weight_rom[6260] = 6;
        weight_rom[6261] = -19;
        weight_rom[6262] = -19;
        weight_rom[6263] = -13;
        weight_rom[6264] = -14;
        weight_rom[6265] = -13;
        weight_rom[6266] = -4;
        weight_rom[6267] = -2;
        weight_rom[6268] = -4;
        weight_rom[6269] = -2;
        weight_rom[6270] = -4;
        weight_rom[6271] = -1;
        weight_rom[6272] = -4;
        weight_rom[6273] = 4;
        weight_rom[6274] = 0;
        weight_rom[6275] = 4;
        weight_rom[6276] = -1;
        weight_rom[6277] = -4;
        weight_rom[6278] = -4;
        weight_rom[6279] = 4;
        weight_rom[6280] = -1;
        weight_rom[6281] = 0;
        weight_rom[6282] = 4;
        weight_rom[6283] = 2;
        weight_rom[6284] = 4;
        weight_rom[6285] = 9;
        weight_rom[6286] = 0;
        weight_rom[6287] = 4;
        weight_rom[6288] = -1;
        weight_rom[6289] = -1;
        weight_rom[6290] = -4;
        weight_rom[6291] = -1;
        weight_rom[6292] = -2;
        weight_rom[6293] = -1;
        weight_rom[6294] = 3;
        weight_rom[6295] = 1;
        weight_rom[6296] = -1;
        weight_rom[6297] = -4;
        weight_rom[6298] = 3;
        weight_rom[6299] = -3;
        weight_rom[6300] = 3;
        weight_rom[6301] = -4;
        weight_rom[6302] = 2;
        weight_rom[6303] = 2;
        weight_rom[6304] = -3;
        weight_rom[6305] = 1;
        weight_rom[6306] = 16;
        weight_rom[6307] = 22;
        weight_rom[6308] = 12;
        weight_rom[6309] = 24;
        weight_rom[6310] = 30;
        weight_rom[6311] = 25;
        weight_rom[6312] = 43;
        weight_rom[6313] = 39;
        weight_rom[6314] = 9;
        weight_rom[6315] = 12;
        weight_rom[6316] = 4;
        weight_rom[6317] = 23;
        weight_rom[6318] = 17;
        weight_rom[6319] = 18;
        weight_rom[6320] = 18;
        weight_rom[6321] = 7;
        weight_rom[6322] = 9;
        weight_rom[6323] = 19;
        weight_rom[6324] = 1;
        weight_rom[6325] = 2;
        weight_rom[6326] = 1;
        weight_rom[6327] = -2;
        weight_rom[6328] = -4;
        weight_rom[6329] = 1;
        weight_rom[6330] = 2;
        weight_rom[6331] = 2;
        weight_rom[6332] = 12;
        weight_rom[6333] = -5;
        weight_rom[6334] = 21;
        weight_rom[6335] = 34;
        weight_rom[6336] = 33;
        weight_rom[6337] = 1;
        weight_rom[6338] = 24;
        weight_rom[6339] = 23;
        weight_rom[6340] = 31;
        weight_rom[6341] = 35;
        weight_rom[6342] = 34;
        weight_rom[6343] = 13;
        weight_rom[6344] = 14;
        weight_rom[6345] = 16;
        weight_rom[6346] = 2;
        weight_rom[6347] = 6;
        weight_rom[6348] = 14;
        weight_rom[6349] = 1;
        weight_rom[6350] = 20;
        weight_rom[6351] = 19;
        weight_rom[6352] = 7;
        weight_rom[6353] = -1;
        weight_rom[6354] = -1;
        weight_rom[6355] = 2;
        weight_rom[6356] = 1;
        weight_rom[6357] = 3;
        weight_rom[6358] = 7;
        weight_rom[6359] = 5;
        weight_rom[6360] = 1;
        weight_rom[6361] = 22;
        weight_rom[6362] = 12;
        weight_rom[6363] = 16;
        weight_rom[6364] = 11;
        weight_rom[6365] = 9;
        weight_rom[6366] = 13;
        weight_rom[6367] = 31;
        weight_rom[6368] = 30;
        weight_rom[6369] = 29;
        weight_rom[6370] = 36;
        weight_rom[6371] = 34;
        weight_rom[6372] = 25;
        weight_rom[6373] = 24;
        weight_rom[6374] = 24;
        weight_rom[6375] = 29;
        weight_rom[6376] = 24;
        weight_rom[6377] = -2;
        weight_rom[6378] = 1;
        weight_rom[6379] = 11;
        weight_rom[6380] = 13;
        weight_rom[6381] = -9;
        weight_rom[6382] = 2;
        weight_rom[6383] = -2;
        weight_rom[6384] = 4;
        weight_rom[6385] = 1;
        weight_rom[6386] = -1;
        weight_rom[6387] = -1;
        weight_rom[6388] = 12;
        weight_rom[6389] = 7;
        weight_rom[6390] = -5;
        weight_rom[6391] = -2;
        weight_rom[6392] = 11;
        weight_rom[6393] = 8;
        weight_rom[6394] = 3;
        weight_rom[6395] = 11;
        weight_rom[6396] = 0;
        weight_rom[6397] = 11;
        weight_rom[6398] = 1;
        weight_rom[6399] = 5;
        weight_rom[6400] = 14;
        weight_rom[6401] = 13;
        weight_rom[6402] = 6;
        weight_rom[6403] = 13;
        weight_rom[6404] = 9;
        weight_rom[6405] = 21;
        weight_rom[6406] = 33;
        weight_rom[6407] = 16;
        weight_rom[6408] = -12;
        weight_rom[6409] = -15;
        weight_rom[6410] = -13;
        weight_rom[6411] = -1;
        weight_rom[6412] = 2;
        weight_rom[6413] = 3;
        weight_rom[6414] = 3;
        weight_rom[6415] = 0;
        weight_rom[6416] = 14;
        weight_rom[6417] = 18;
        weight_rom[6418] = 33;
        weight_rom[6419] = 10;
        weight_rom[6420] = 6;
        weight_rom[6421] = 7;
        weight_rom[6422] = 9;
        weight_rom[6423] = -12;
        weight_rom[6424] = -8;
        weight_rom[6425] = -8;
        weight_rom[6426] = 7;
        weight_rom[6427] = 10;
        weight_rom[6428] = 8;
        weight_rom[6429] = 6;
        weight_rom[6430] = 24;
        weight_rom[6431] = 20;
        weight_rom[6432] = 13;
        weight_rom[6433] = 4;
        weight_rom[6434] = 11;
        weight_rom[6435] = 15;
        weight_rom[6436] = 4;
        weight_rom[6437] = -10;
        weight_rom[6438] = -4;
        weight_rom[6439] = 1;
        weight_rom[6440] = -4;
        weight_rom[6441] = 0;
        weight_rom[6442] = 12;
        weight_rom[6443] = 5;
        weight_rom[6444] = 30;
        weight_rom[6445] = 9;
        weight_rom[6446] = 8;
        weight_rom[6447] = -9;
        weight_rom[6448] = 12;
        weight_rom[6449] = 3;
        weight_rom[6450] = -5;
        weight_rom[6451] = -17;
        weight_rom[6452] = -7;
        weight_rom[6453] = -11;
        weight_rom[6454] = -15;
        weight_rom[6455] = -13;
        weight_rom[6456] = -15;
        weight_rom[6457] = -10;
        weight_rom[6458] = -2;
        weight_rom[6459] = -8;
        weight_rom[6460] = 5;
        weight_rom[6461] = 13;
        weight_rom[6462] = 13;
        weight_rom[6463] = 34;
        weight_rom[6464] = 10;
        weight_rom[6465] = 4;
        weight_rom[6466] = 2;
        weight_rom[6467] = -14;
        weight_rom[6468] = 2;
        weight_rom[6469] = 2;
        weight_rom[6470] = -7;
        weight_rom[6471] = 14;
        weight_rom[6472] = 16;
        weight_rom[6473] = 18;
        weight_rom[6474] = 6;
        weight_rom[6475] = 23;
        weight_rom[6476] = -13;
        weight_rom[6477] = -14;
        weight_rom[6478] = -15;
        weight_rom[6479] = -11;
        weight_rom[6480] = -11;
        weight_rom[6481] = -18;
        weight_rom[6482] = -16;
        weight_rom[6483] = -21;
        weight_rom[6484] = -28;
        weight_rom[6485] = -12;
        weight_rom[6486] = -6;
        weight_rom[6487] = -5;
        weight_rom[6488] = -19;
        weight_rom[6489] = -4;
        weight_rom[6490] = 5;
        weight_rom[6491] = 11;
        weight_rom[6492] = 29;
        weight_rom[6493] = 10;
        weight_rom[6494] = 8;
        weight_rom[6495] = 17;
        weight_rom[6496] = 16;
        weight_rom[6497] = 18;
        weight_rom[6498] = 18;
        weight_rom[6499] = 18;
        weight_rom[6500] = 18;
        weight_rom[6501] = 18;
        weight_rom[6502] = 3;
        weight_rom[6503] = -3;
        weight_rom[6504] = -8;
        weight_rom[6505] = 0;
        weight_rom[6506] = -9;
        weight_rom[6507] = -5;
        weight_rom[6508] = 10;
        weight_rom[6509] = 4;
        weight_rom[6510] = -10;
        weight_rom[6511] = -11;
        weight_rom[6512] = -15;
        weight_rom[6513] = -15;
        weight_rom[6514] = -8;
        weight_rom[6515] = -15;
        weight_rom[6516] = -1;
        weight_rom[6517] = -5;
        weight_rom[6518] = 1;
        weight_rom[6519] = 3;
        weight_rom[6520] = 12;
        weight_rom[6521] = 9;
        weight_rom[6522] = -20;
        weight_rom[6523] = -14;
        weight_rom[6524] = 10;
        weight_rom[6525] = 21;
        weight_rom[6526] = 18;
        weight_rom[6527] = 18;
        weight_rom[6528] = 22;
        weight_rom[6529] = 2;
        weight_rom[6530] = -8;
        weight_rom[6531] = -1;
        weight_rom[6532] = -7;
        weight_rom[6533] = -7;
        weight_rom[6534] = -1;
        weight_rom[6535] = 11;
        weight_rom[6536] = 16;
        weight_rom[6537] = 25;
        weight_rom[6538] = 10;
        weight_rom[6539] = -8;
        weight_rom[6540] = -14;
        weight_rom[6541] = -15;
        weight_rom[6542] = -4;
        weight_rom[6543] = -7;
        weight_rom[6544] = -6;
        weight_rom[6545] = 9;
        weight_rom[6546] = 1;
        weight_rom[6547] = 4;
        weight_rom[6548] = 9;
        weight_rom[6549] = 5;
        weight_rom[6550] = -4;
        weight_rom[6551] = 2;
        weight_rom[6552] = 17;
        weight_rom[6553] = 20;
        weight_rom[6554] = 23;
        weight_rom[6555] = 19;
        weight_rom[6556] = 4;
        weight_rom[6557] = 0;
        weight_rom[6558] = -11;
        weight_rom[6559] = -5;
        weight_rom[6560] = -5;
        weight_rom[6561] = 2;
        weight_rom[6562] = 9;
        weight_rom[6563] = 26;
        weight_rom[6564] = 36;
        weight_rom[6565] = 38;
        weight_rom[6566] = 6;
        weight_rom[6567] = -9;
        weight_rom[6568] = -16;
        weight_rom[6569] = -3;
        weight_rom[6570] = -4;
        weight_rom[6571] = 1;
        weight_rom[6572] = 9;
        weight_rom[6573] = 10;
        weight_rom[6574] = 12;
        weight_rom[6575] = -2;
        weight_rom[6576] = 6;
        weight_rom[6577] = 33;
        weight_rom[6578] = -23;
        weight_rom[6579] = -12;
        weight_rom[6580] = 21;
        weight_rom[6581] = 25;
        weight_rom[6582] = 46;
        weight_rom[6583] = 22;
        weight_rom[6584] = 15;
        weight_rom[6585] = -7;
        weight_rom[6586] = -6;
        weight_rom[6587] = 13;
        weight_rom[6588] = 10;
        weight_rom[6589] = 23;
        weight_rom[6590] = 37;
        weight_rom[6591] = 50;
        weight_rom[6592] = 55;
        weight_rom[6593] = 24;
        weight_rom[6594] = -5;
        weight_rom[6595] = -17;
        weight_rom[6596] = -4;
        weight_rom[6597] = -2;
        weight_rom[6598] = 3;
        weight_rom[6599] = -2;
        weight_rom[6600] = -4;
        weight_rom[6601] = 3;
        weight_rom[6602] = 10;
        weight_rom[6603] = 6;
        weight_rom[6604] = 2;
        weight_rom[6605] = -1;
        weight_rom[6606] = -6;
        weight_rom[6607] = 16;
        weight_rom[6608] = 8;
        weight_rom[6609] = 20;
        weight_rom[6610] = 33;
        weight_rom[6611] = 29;
        weight_rom[6612] = -4;
        weight_rom[6613] = -8;
        weight_rom[6614] = 10;
        weight_rom[6615] = 32;
        weight_rom[6616] = 37;
        weight_rom[6617] = 50;
        weight_rom[6618] = 55;
        weight_rom[6619] = 54;
        weight_rom[6620] = 26;
        weight_rom[6621] = 2;
        weight_rom[6622] = -20;
        weight_rom[6623] = -14;
        weight_rom[6624] = 3;
        weight_rom[6625] = 9;
        weight_rom[6626] = 3;
        weight_rom[6627] = -12;
        weight_rom[6628] = -16;
        weight_rom[6629] = 3;
        weight_rom[6630] = 15;
        weight_rom[6631] = 12;
        weight_rom[6632] = 14;
        weight_rom[6633] = -6;
        weight_rom[6634] = -19;
        weight_rom[6635] = 13;
        weight_rom[6636] = -1;
        weight_rom[6637] = 1;
        weight_rom[6638] = 39;
        weight_rom[6639] = 4;
        weight_rom[6640] = 7;
        weight_rom[6641] = 24;
        weight_rom[6642] = 41;
        weight_rom[6643] = 48;
        weight_rom[6644] = 39;
        weight_rom[6645] = 50;
        weight_rom[6646] = 43;
        weight_rom[6647] = 21;
        weight_rom[6648] = -20;
        weight_rom[6649] = -29;
        weight_rom[6650] = -20;
        weight_rom[6651] = -15;
        weight_rom[6652] = 2;
        weight_rom[6653] = 7;
        weight_rom[6654] = 0;
        weight_rom[6655] = -7;
        weight_rom[6656] = -5;
        weight_rom[6657] = 13;
        weight_rom[6658] = 13;
        weight_rom[6659] = 31;
        weight_rom[6660] = 10;
        weight_rom[6661] = -8;
        weight_rom[6662] = -22;
        weight_rom[6663] = -20;
        weight_rom[6664] = -1;
        weight_rom[6665] = 4;
        weight_rom[6666] = 20;
        weight_rom[6667] = 16;
        weight_rom[6668] = 12;
        weight_rom[6669] = 39;
        weight_rom[6670] = 36;
        weight_rom[6671] = 35;
        weight_rom[6672] = 34;
        weight_rom[6673] = 25;
        weight_rom[6674] = 7;
        weight_rom[6675] = -16;
        weight_rom[6676] = -34;
        weight_rom[6677] = -46;
        weight_rom[6678] = -20;
        weight_rom[6679] = -11;
        weight_rom[6680] = -3;
        weight_rom[6681] = 0;
        weight_rom[6682] = -6;
        weight_rom[6683] = -8;
        weight_rom[6684] = 9;
        weight_rom[6685] = 15;
        weight_rom[6686] = 33;
        weight_rom[6687] = 44;
        weight_rom[6688] = 30;
        weight_rom[6689] = -23;
        weight_rom[6690] = -27;
        weight_rom[6691] = -2;
        weight_rom[6692] = 3;
        weight_rom[6693] = 1;
        weight_rom[6694] = 28;
        weight_rom[6695] = 7;
        weight_rom[6696] = 2;
        weight_rom[6697] = 33;
        weight_rom[6698] = 28;
        weight_rom[6699] = 26;
        weight_rom[6700] = 12;
        weight_rom[6701] = 7;
        weight_rom[6702] = -10;
        weight_rom[6703] = -26;
        weight_rom[6704] = -26;
        weight_rom[6705] = -41;
        weight_rom[6706] = -23;
        weight_rom[6707] = -5;
        weight_rom[6708] = -12;
        weight_rom[6709] = 1;
        weight_rom[6710] = -3;
        weight_rom[6711] = -3;
        weight_rom[6712] = 15;
        weight_rom[6713] = 21;
        weight_rom[6714] = 36;
        weight_rom[6715] = 44;
        weight_rom[6716] = 2;
        weight_rom[6717] = -26;
        weight_rom[6718] = -29;
        weight_rom[6719] = -5;
        weight_rom[6720] = 1;
        weight_rom[6721] = 2;
        weight_rom[6722] = 17;
        weight_rom[6723] = -10;
        weight_rom[6724] = -11;
        weight_rom[6725] = 6;
        weight_rom[6726] = 7;
        weight_rom[6727] = 17;
        weight_rom[6728] = 15;
        weight_rom[6729] = -9;
        weight_rom[6730] = -19;
        weight_rom[6731] = -25;
        weight_rom[6732] = -41;
        weight_rom[6733] = -38;
        weight_rom[6734] = -19;
        weight_rom[6735] = -2;
        weight_rom[6736] = -8;
        weight_rom[6737] = -10;
        weight_rom[6738] = -9;
        weight_rom[6739] = 11;
        weight_rom[6740] = 9;
        weight_rom[6741] = 22;
        weight_rom[6742] = 16;
        weight_rom[6743] = 19;
        weight_rom[6744] = 2;
        weight_rom[6745] = -42;
        weight_rom[6746] = -33;
        weight_rom[6747] = -20;
        weight_rom[6748] = 4;
        weight_rom[6749] = 8;
        weight_rom[6750] = 2;
        weight_rom[6751] = -8;
        weight_rom[6752] = -3;
        weight_rom[6753] = 1;
        weight_rom[6754] = 2;
        weight_rom[6755] = 3;
        weight_rom[6756] = 3;
        weight_rom[6757] = -5;
        weight_rom[6758] = -11;
        weight_rom[6759] = -20;
        weight_rom[6760] = -34;
        weight_rom[6761] = -43;
        weight_rom[6762] = -10;
        weight_rom[6763] = -1;
        weight_rom[6764] = -5;
        weight_rom[6765] = 0;
        weight_rom[6766] = 0;
        weight_rom[6767] = 1;
        weight_rom[6768] = 10;
        weight_rom[6769] = 24;
        weight_rom[6770] = 19;
        weight_rom[6771] = 17;
        weight_rom[6772] = -14;
        weight_rom[6773] = -31;
        weight_rom[6774] = -30;
        weight_rom[6775] = -3;
        weight_rom[6776] = -1;
        weight_rom[6777] = 7;
        weight_rom[6778] = 4;
        weight_rom[6779] = 18;
        weight_rom[6780] = -4;
        weight_rom[6781] = -19;
        weight_rom[6782] = -8;
        weight_rom[6783] = -1;
        weight_rom[6784] = 6;
        weight_rom[6785] = 12;
        weight_rom[6786] = -2;
        weight_rom[6787] = -5;
        weight_rom[6788] = -35;
        weight_rom[6789] = -42;
        weight_rom[6790] = -11;
        weight_rom[6791] = -2;
        weight_rom[6792] = 1;
        weight_rom[6793] = 8;
        weight_rom[6794] = 4;
        weight_rom[6795] = 12;
        weight_rom[6796] = 14;
        weight_rom[6797] = 30;
        weight_rom[6798] = 9;
        weight_rom[6799] = -9;
        weight_rom[6800] = -22;
        weight_rom[6801] = -15;
        weight_rom[6802] = -9;
        weight_rom[6803] = -14;
        weight_rom[6804] = 3;
        weight_rom[6805] = 8;
        weight_rom[6806] = -7;
        weight_rom[6807] = 18;
        weight_rom[6808] = -14;
        weight_rom[6809] = -18;
        weight_rom[6810] = -18;
        weight_rom[6811] = -16;
        weight_rom[6812] = -1;
        weight_rom[6813] = 8;
        weight_rom[6814] = 1;
        weight_rom[6815] = 0;
        weight_rom[6816] = -6;
        weight_rom[6817] = -18;
        weight_rom[6818] = 11;
        weight_rom[6819] = 9;
        weight_rom[6820] = 24;
        weight_rom[6821] = 13;
        weight_rom[6822] = 15;
        weight_rom[6823] = 12;
        weight_rom[6824] = 19;
        weight_rom[6825] = 13;
        weight_rom[6826] = -4;
        weight_rom[6827] = -18;
        weight_rom[6828] = 1;
        weight_rom[6829] = -16;
        weight_rom[6830] = -16;
        weight_rom[6831] = -9;
        weight_rom[6832] = -2;
        weight_rom[6833] = 14;
        weight_rom[6834] = -4;
        weight_rom[6835] = -9;
        weight_rom[6836] = -26;
        weight_rom[6837] = -31;
        weight_rom[6838] = -22;
        weight_rom[6839] = -16;
        weight_rom[6840] = -1;
        weight_rom[6841] = 8;
        weight_rom[6842] = 17;
        weight_rom[6843] = 16;
        weight_rom[6844] = 11;
        weight_rom[6845] = 3;
        weight_rom[6846] = 17;
        weight_rom[6847] = 20;
        weight_rom[6848] = 20;
        weight_rom[6849] = 25;
        weight_rom[6850] = 19;
        weight_rom[6851] = 18;
        weight_rom[6852] = 10;
        weight_rom[6853] = -7;
        weight_rom[6854] = -22;
        weight_rom[6855] = -20;
        weight_rom[6856] = -9;
        weight_rom[6857] = -30;
        weight_rom[6858] = 1;
        weight_rom[6859] = 1;
        weight_rom[6860] = -2;
        weight_rom[6861] = 0;
        weight_rom[6862] = -7;
        weight_rom[6863] = -8;
        weight_rom[6864] = -33;
        weight_rom[6865] = -26;
        weight_rom[6866] = -36;
        weight_rom[6867] = -24;
        weight_rom[6868] = -12;
        weight_rom[6869] = -15;
        weight_rom[6870] = 1;
        weight_rom[6871] = 9;
        weight_rom[6872] = 10;
        weight_rom[6873] = 6;
        weight_rom[6874] = 16;
        weight_rom[6875] = 26;
        weight_rom[6876] = 20;
        weight_rom[6877] = 20;
        weight_rom[6878] = 23;
        weight_rom[6879] = 6;
        weight_rom[6880] = 0;
        weight_rom[6881] = -10;
        weight_rom[6882] = -16;
        weight_rom[6883] = -33;
        weight_rom[6884] = -25;
        weight_rom[6885] = -19;
        weight_rom[6886] = 8;
        weight_rom[6887] = 0;
        weight_rom[6888] = 0;
        weight_rom[6889] = -3;
        weight_rom[6890] = -1;
        weight_rom[6891] = -6;
        weight_rom[6892] = -13;
        weight_rom[6893] = -15;
        weight_rom[6894] = -27;
        weight_rom[6895] = -25;
        weight_rom[6896] = -15;
        weight_rom[6897] = -6;
        weight_rom[6898] = -2;
        weight_rom[6899] = 3;
        weight_rom[6900] = 3;
        weight_rom[6901] = 12;
        weight_rom[6902] = 9;
        weight_rom[6903] = 15;
        weight_rom[6904] = 11;
        weight_rom[6905] = 22;
        weight_rom[6906] = 11;
        weight_rom[6907] = 22;
        weight_rom[6908] = -2;
        weight_rom[6909] = -5;
        weight_rom[6910] = -11;
        weight_rom[6911] = -28;
        weight_rom[6912] = -31;
        weight_rom[6913] = -14;
        weight_rom[6914] = 2;
        weight_rom[6915] = -1;
        weight_rom[6916] = 1;
        weight_rom[6917] = 2;
        weight_rom[6918] = 9;
        weight_rom[6919] = 18;
        weight_rom[6920] = 10;
        weight_rom[6921] = 1;
        weight_rom[6922] = 3;
        weight_rom[6923] = 5;
        weight_rom[6924] = -15;
        weight_rom[6925] = 0;
        weight_rom[6926] = 7;
        weight_rom[6927] = 1;
        weight_rom[6928] = -4;
        weight_rom[6929] = -8;
        weight_rom[6930] = 9;
        weight_rom[6931] = 19;
        weight_rom[6932] = 8;
        weight_rom[6933] = 9;
        weight_rom[6934] = 17;
        weight_rom[6935] = 2;
        weight_rom[6936] = -2;
        weight_rom[6937] = -4;
        weight_rom[6938] = -49;
        weight_rom[6939] = -52;
        weight_rom[6940] = -39;
        weight_rom[6941] = -19;
        weight_rom[6942] = 2;
        weight_rom[6943] = -1;
        weight_rom[6944] = -2;
        weight_rom[6945] = 2;
        weight_rom[6946] = 5;
        weight_rom[6947] = 12;
        weight_rom[6948] = 29;
        weight_rom[6949] = 28;
        weight_rom[6950] = 8;
        weight_rom[6951] = 12;
        weight_rom[6952] = 9;
        weight_rom[6953] = 5;
        weight_rom[6954] = 14;
        weight_rom[6955] = 6;
        weight_rom[6956] = 2;
        weight_rom[6957] = 7;
        weight_rom[6958] = 4;
        weight_rom[6959] = 3;
        weight_rom[6960] = 15;
        weight_rom[6961] = 16;
        weight_rom[6962] = -1;
        weight_rom[6963] = 4;
        weight_rom[6964] = -14;
        weight_rom[6965] = -22;
        weight_rom[6966] = -15;
        weight_rom[6967] = -18;
        weight_rom[6968] = -14;
        weight_rom[6969] = -4;
        weight_rom[6970] = 3;
        weight_rom[6971] = 4;
        weight_rom[6972] = -3;
        weight_rom[6973] = -4;
        weight_rom[6974] = -1;
        weight_rom[6975] = -19;
        weight_rom[6976] = 15;
        weight_rom[6977] = 8;
        weight_rom[6978] = 24;
        weight_rom[6979] = 7;
        weight_rom[6980] = 17;
        weight_rom[6981] = 3;
        weight_rom[6982] = 1;
        weight_rom[6983] = 7;
        weight_rom[6984] = 4;
        weight_rom[6985] = -6;
        weight_rom[6986] = -10;
        weight_rom[6987] = -4;
        weight_rom[6988] = 0;
        weight_rom[6989] = -5;
        weight_rom[6990] = 8;
        weight_rom[6991] = -10;
        weight_rom[6992] = -16;
        weight_rom[6993] = -6;
        weight_rom[6994] = -2;
        weight_rom[6995] = 6;
        weight_rom[6996] = -11;
        weight_rom[6997] = 4;
        weight_rom[6998] = 3;
        weight_rom[6999] = -2;
        weight_rom[7000] = 2;
        weight_rom[7001] = 1;
        weight_rom[7002] = 1;
        weight_rom[7003] = 2;
        weight_rom[7004] = -7;
        weight_rom[7005] = -24;
        weight_rom[7006] = -22;
        weight_rom[7007] = -13;
        weight_rom[7008] = -2;
        weight_rom[7009] = -7;
        weight_rom[7010] = -15;
        weight_rom[7011] = -8;
        weight_rom[7012] = -16;
        weight_rom[7013] = -12;
        weight_rom[7014] = -21;
        weight_rom[7015] = 1;
        weight_rom[7016] = 0;
        weight_rom[7017] = -4;
        weight_rom[7018] = -13;
        weight_rom[7019] = 8;
        weight_rom[7020] = -9;
        weight_rom[7021] = -12;
        weight_rom[7022] = -3;
        weight_rom[7023] = -12;
        weight_rom[7024] = 4;
        weight_rom[7025] = -4;
        weight_rom[7026] = 1;
        weight_rom[7027] = -1;
        weight_rom[7028] = -1;
        weight_rom[7029] = -2;
        weight_rom[7030] = -3;
        weight_rom[7031] = 4;
        weight_rom[7032] = -2;
        weight_rom[7033] = 18;
        weight_rom[7034] = 20;
        weight_rom[7035] = -8;
        weight_rom[7036] = -8;
        weight_rom[7037] = 1;
        weight_rom[7038] = 2;
        weight_rom[7039] = -6;
        weight_rom[7040] = 4;
        weight_rom[7041] = 47;
        weight_rom[7042] = 6;
        weight_rom[7043] = 4;
        weight_rom[7044] = 10;
        weight_rom[7045] = 43;
        weight_rom[7046] = 15;
        weight_rom[7047] = -5;
        weight_rom[7048] = 8;
        weight_rom[7049] = 6;
        weight_rom[7050] = 19;
        weight_rom[7051] = -4;
        weight_rom[7052] = 2;
        weight_rom[7053] = 2;
        weight_rom[7054] = 1;
        weight_rom[7055] = 4;
        weight_rom[7056] = 2;
        weight_rom[7057] = 4;
        weight_rom[7058] = 3;
        weight_rom[7059] = 3;
        weight_rom[7060] = 3;
        weight_rom[7061] = 4;
        weight_rom[7062] = -1;
        weight_rom[7063] = 3;
        weight_rom[7064] = 1;
        weight_rom[7065] = 4;
        weight_rom[7066] = 0;
        weight_rom[7067] = -2;
        weight_rom[7068] = 0;
        weight_rom[7069] = -3;
        weight_rom[7070] = 4;
        weight_rom[7071] = -1;
        weight_rom[7072] = -3;
        weight_rom[7073] = -3;
        weight_rom[7074] = -3;
        weight_rom[7075] = -2;
        weight_rom[7076] = -3;
        weight_rom[7077] = 0;
        weight_rom[7078] = -3;
        weight_rom[7079] = -3;
        weight_rom[7080] = 4;
        weight_rom[7081] = 4;
        weight_rom[7082] = -4;
        weight_rom[7083] = -1;
        weight_rom[7084] = 4;
        weight_rom[7085] = 1;
        weight_rom[7086] = 4;
        weight_rom[7087] = 3;
        weight_rom[7088] = -4;
        weight_rom[7089] = 2;
        weight_rom[7090] = -14;
        weight_rom[7091] = -20;
        weight_rom[7092] = -7;
        weight_rom[7093] = -7;
        weight_rom[7094] = -4;
        weight_rom[7095] = -10;
        weight_rom[7096] = -17;
        weight_rom[7097] = -7;
        weight_rom[7098] = 4;
        weight_rom[7099] = -3;
        weight_rom[7100] = -8;
        weight_rom[7101] = 9;
        weight_rom[7102] = 4;
        weight_rom[7103] = 7;
        weight_rom[7104] = -1;
        weight_rom[7105] = -6;
        weight_rom[7106] = -11;
        weight_rom[7107] = -11;
        weight_rom[7108] = -1;
        weight_rom[7109] = 1;
        weight_rom[7110] = 0;
        weight_rom[7111] = -3;
        weight_rom[7112] = 1;
        weight_rom[7113] = 1;
        weight_rom[7114] = 2;
        weight_rom[7115] = -1;
        weight_rom[7116] = -2;
        weight_rom[7117] = -1;
        weight_rom[7118] = -7;
        weight_rom[7119] = -12;
        weight_rom[7120] = 5;
        weight_rom[7121] = 38;
        weight_rom[7122] = 29;
        weight_rom[7123] = 41;
        weight_rom[7124] = 16;
        weight_rom[7125] = 1;
        weight_rom[7126] = 18;
        weight_rom[7127] = 23;
        weight_rom[7128] = 16;
        weight_rom[7129] = 26;
        weight_rom[7130] = 12;
        weight_rom[7131] = 23;
        weight_rom[7132] = 28;
        weight_rom[7133] = 15;
        weight_rom[7134] = 19;
        weight_rom[7135] = 21;
        weight_rom[7136] = 27;
        weight_rom[7137] = 16;
        weight_rom[7138] = -2;
        weight_rom[7139] = -4;
        weight_rom[7140] = 4;
        weight_rom[7141] = 2;
        weight_rom[7142] = 2;
        weight_rom[7143] = -3;
        weight_rom[7144] = -3;
        weight_rom[7145] = 1;
        weight_rom[7146] = 25;
        weight_rom[7147] = 9;
        weight_rom[7148] = -1;
        weight_rom[7149] = 15;
        weight_rom[7150] = 5;
        weight_rom[7151] = 7;
        weight_rom[7152] = 0;
        weight_rom[7153] = -8;
        weight_rom[7154] = -8;
        weight_rom[7155] = -4;
        weight_rom[7156] = -7;
        weight_rom[7157] = 11;
        weight_rom[7158] = 16;
        weight_rom[7159] = 23;
        weight_rom[7160] = 15;
        weight_rom[7161] = 21;
        weight_rom[7162] = 17;
        weight_rom[7163] = 7;
        weight_rom[7164] = 18;
        weight_rom[7165] = 4;
        weight_rom[7166] = -3;
        weight_rom[7167] = 4;
        weight_rom[7168] = 2;
        weight_rom[7169] = -2;
        weight_rom[7170] = -9;
        weight_rom[7171] = -4;
        weight_rom[7172] = 7;
        weight_rom[7173] = 8;
        weight_rom[7174] = 12;
        weight_rom[7175] = 8;
        weight_rom[7176] = 10;
        weight_rom[7177] = -15;
        weight_rom[7178] = -14;
        weight_rom[7179] = -6;
        weight_rom[7180] = -8;
        weight_rom[7181] = -26;
        weight_rom[7182] = -32;
        weight_rom[7183] = -35;
        weight_rom[7184] = -29;
        weight_rom[7185] = -8;
        weight_rom[7186] = -16;
        weight_rom[7187] = -15;
        weight_rom[7188] = -11;
        weight_rom[7189] = -6;
        weight_rom[7190] = 13;
        weight_rom[7191] = 4;
        weight_rom[7192] = -5;
        weight_rom[7193] = 3;
        weight_rom[7194] = -8;
        weight_rom[7195] = 2;
        weight_rom[7196] = 1;
        weight_rom[7197] = -5;
        weight_rom[7198] = 1;
        weight_rom[7199] = 3;
        weight_rom[7200] = 16;
        weight_rom[7201] = 2;
        weight_rom[7202] = 9;
        weight_rom[7203] = -4;
        weight_rom[7204] = 15;
        weight_rom[7205] = 20;
        weight_rom[7206] = -2;
        weight_rom[7207] = -10;
        weight_rom[7208] = -23;
        weight_rom[7209] = -16;
        weight_rom[7210] = -14;
        weight_rom[7211] = -25;
        weight_rom[7212] = -20;
        weight_rom[7213] = -11;
        weight_rom[7214] = -6;
        weight_rom[7215] = -16;
        weight_rom[7216] = -19;
        weight_rom[7217] = -22;
        weight_rom[7218] = -17;
        weight_rom[7219] = -3;
        weight_rom[7220] = 5;
        weight_rom[7221] = -13;
        weight_rom[7222] = -25;
        weight_rom[7223] = 4;
        weight_rom[7224] = 1;
        weight_rom[7225] = -2;
        weight_rom[7226] = -12;
        weight_rom[7227] = -5;
        weight_rom[7228] = 23;
        weight_rom[7229] = 12;
        weight_rom[7230] = 13;
        weight_rom[7231] = 21;
        weight_rom[7232] = 13;
        weight_rom[7233] = 5;
        weight_rom[7234] = -5;
        weight_rom[7235] = -10;
        weight_rom[7236] = -15;
        weight_rom[7237] = -18;
        weight_rom[7238] = -2;
        weight_rom[7239] = 0;
        weight_rom[7240] = -2;
        weight_rom[7241] = 5;
        weight_rom[7242] = -14;
        weight_rom[7243] = -23;
        weight_rom[7244] = -28;
        weight_rom[7245] = -22;
        weight_rom[7246] = -22;
        weight_rom[7247] = -14;
        weight_rom[7248] = -26;
        weight_rom[7249] = -12;
        weight_rom[7250] = -2;
        weight_rom[7251] = -8;
        weight_rom[7252] = 1;
        weight_rom[7253] = -18;
        weight_rom[7254] = 30;
        weight_rom[7255] = 2;
        weight_rom[7256] = 5;
        weight_rom[7257] = 7;
        weight_rom[7258] = 22;
        weight_rom[7259] = 12;
        weight_rom[7260] = -9;
        weight_rom[7261] = 7;
        weight_rom[7262] = -1;
        weight_rom[7263] = -8;
        weight_rom[7264] = -4;
        weight_rom[7265] = 2;
        weight_rom[7266] = 10;
        weight_rom[7267] = 8;
        weight_rom[7268] = 11;
        weight_rom[7269] = 3;
        weight_rom[7270] = -15;
        weight_rom[7271] = -22;
        weight_rom[7272] = -11;
        weight_rom[7273] = -17;
        weight_rom[7274] = -12;
        weight_rom[7275] = -34;
        weight_rom[7276] = -14;
        weight_rom[7277] = -5;
        weight_rom[7278] = 7;
        weight_rom[7279] = -9;
        weight_rom[7280] = 13;
        weight_rom[7281] = 9;
        weight_rom[7282] = 20;
        weight_rom[7283] = -1;
        weight_rom[7284] = 8;
        weight_rom[7285] = 16;
        weight_rom[7286] = 5;
        weight_rom[7287] = -10;
        weight_rom[7288] = 8;
        weight_rom[7289] = 2;
        weight_rom[7290] = -3;
        weight_rom[7291] = 1;
        weight_rom[7292] = -3;
        weight_rom[7293] = -4;
        weight_rom[7294] = -1;
        weight_rom[7295] = 0;
        weight_rom[7296] = -13;
        weight_rom[7297] = -7;
        weight_rom[7298] = -23;
        weight_rom[7299] = -26;
        weight_rom[7300] = -23;
        weight_rom[7301] = -15;
        weight_rom[7302] = -19;
        weight_rom[7303] = -27;
        weight_rom[7304] = -19;
        weight_rom[7305] = -15;
        weight_rom[7306] = -27;
        weight_rom[7307] = -15;
        weight_rom[7308] = 8;
        weight_rom[7309] = 11;
        weight_rom[7310] = 14;
        weight_rom[7311] = 2;
        weight_rom[7312] = 10;
        weight_rom[7313] = 13;
        weight_rom[7314] = 10;
        weight_rom[7315] = 4;
        weight_rom[7316] = -6;
        weight_rom[7317] = -8;
        weight_rom[7318] = 4;
        weight_rom[7319] = 8;
        weight_rom[7320] = 16;
        weight_rom[7321] = 7;
        weight_rom[7322] = 1;
        weight_rom[7323] = -4;
        weight_rom[7324] = -1;
        weight_rom[7325] = -4;
        weight_rom[7326] = -12;
        weight_rom[7327] = -11;
        weight_rom[7328] = -15;
        weight_rom[7329] = -17;
        weight_rom[7330] = -28;
        weight_rom[7331] = -31;
        weight_rom[7332] = -35;
        weight_rom[7333] = -46;
        weight_rom[7334] = -15;
        weight_rom[7335] = 9;
        weight_rom[7336] = 17;
        weight_rom[7337] = 21;
        weight_rom[7338] = 4;
        weight_rom[7339] = -4;
        weight_rom[7340] = -23;
        weight_rom[7341] = 9;
        weight_rom[7342] = 8;
        weight_rom[7343] = -4;
        weight_rom[7344] = 4;
        weight_rom[7345] = 6;
        weight_rom[7346] = 11;
        weight_rom[7347] = 13;
        weight_rom[7348] = 21;
        weight_rom[7349] = 6;
        weight_rom[7350] = -24;
        weight_rom[7351] = -15;
        weight_rom[7352] = -10;
        weight_rom[7353] = -1;
        weight_rom[7354] = -3;
        weight_rom[7355] = -4;
        weight_rom[7356] = -13;
        weight_rom[7357] = -21;
        weight_rom[7358] = -24;
        weight_rom[7359] = -52;
        weight_rom[7360] = -59;
        weight_rom[7361] = -32;
        weight_rom[7362] = -29;
        weight_rom[7363] = -20;
        weight_rom[7364] = 14;
        weight_rom[7365] = 15;
        weight_rom[7366] = 13;
        weight_rom[7367] = 7;
        weight_rom[7368] = -10;
        weight_rom[7369] = 0;
        weight_rom[7370] = 4;
        weight_rom[7371] = -1;
        weight_rom[7372] = -1;
        weight_rom[7373] = 9;
        weight_rom[7374] = 9;
        weight_rom[7375] = 19;
        weight_rom[7376] = 25;
        weight_rom[7377] = -22;
        weight_rom[7378] = -31;
        weight_rom[7379] = -15;
        weight_rom[7380] = 12;
        weight_rom[7381] = 5;
        weight_rom[7382] = 3;
        weight_rom[7383] = 11;
        weight_rom[7384] = 15;
        weight_rom[7385] = -3;
        weight_rom[7386] = -23;
        weight_rom[7387] = -49;
        weight_rom[7388] = -54;
        weight_rom[7389] = -41;
        weight_rom[7390] = -43;
        weight_rom[7391] = 12;
        weight_rom[7392] = 14;
        weight_rom[7393] = 10;
        weight_rom[7394] = 17;
        weight_rom[7395] = -6;
        weight_rom[7396] = -8;
        weight_rom[7397] = -3;
        weight_rom[7398] = -5;
        weight_rom[7399] = -2;
        weight_rom[7400] = 4;
        weight_rom[7401] = -2;
        weight_rom[7402] = 7;
        weight_rom[7403] = 19;
        weight_rom[7404] = 11;
        weight_rom[7405] = -16;
        weight_rom[7406] = -17;
        weight_rom[7407] = -7;
        weight_rom[7408] = 22;
        weight_rom[7409] = 18;
        weight_rom[7410] = 13;
        weight_rom[7411] = 20;
        weight_rom[7412] = 12;
        weight_rom[7413] = 1;
        weight_rom[7414] = 3;
        weight_rom[7415] = -21;
        weight_rom[7416] = -32;
        weight_rom[7417] = -19;
        weight_rom[7418] = -26;
        weight_rom[7419] = 18;
        weight_rom[7420] = -5;
        weight_rom[7421] = 3;
        weight_rom[7422] = -4;
        weight_rom[7423] = -11;
        weight_rom[7424] = 12;
        weight_rom[7425] = 3;
        weight_rom[7426] = -1;
        weight_rom[7427] = 1;
        weight_rom[7428] = 10;
        weight_rom[7429] = 5;
        weight_rom[7430] = 22;
        weight_rom[7431] = 20;
        weight_rom[7432] = -7;
        weight_rom[7433] = -6;
        weight_rom[7434] = -4;
        weight_rom[7435] = 11;
        weight_rom[7436] = 33;
        weight_rom[7437] = 32;
        weight_rom[7438] = 30;
        weight_rom[7439] = 24;
        weight_rom[7440] = 26;
        weight_rom[7441] = 18;
        weight_rom[7442] = -7;
        weight_rom[7443] = -11;
        weight_rom[7444] = 0;
        weight_rom[7445] = -3;
        weight_rom[7446] = 2;
        weight_rom[7447] = 13;
        weight_rom[7448] = 0;
        weight_rom[7449] = -7;
        weight_rom[7450] = 14;
        weight_rom[7451] = 1;
        weight_rom[7452] = 20;
        weight_rom[7453] = 6;
        weight_rom[7454] = 5;
        weight_rom[7455] = 18;
        weight_rom[7456] = 10;
        weight_rom[7457] = 22;
        weight_rom[7458] = 20;
        weight_rom[7459] = 28;
        weight_rom[7460] = 7;
        weight_rom[7461] = -9;
        weight_rom[7462] = -1;
        weight_rom[7463] = 15;
        weight_rom[7464] = 42;
        weight_rom[7465] = 41;
        weight_rom[7466] = 44;
        weight_rom[7467] = 43;
        weight_rom[7468] = 36;
        weight_rom[7469] = 6;
        weight_rom[7470] = 17;
        weight_rom[7471] = 6;
        weight_rom[7472] = -28;
        weight_rom[7473] = 25;
        weight_rom[7474] = 21;
        weight_rom[7475] = 4;
        weight_rom[7476] = -1;
        weight_rom[7477] = -9;
        weight_rom[7478] = -2;
        weight_rom[7479] = 16;
        weight_rom[7480] = 1;
        weight_rom[7481] = 0;
        weight_rom[7482] = 27;
        weight_rom[7483] = 10;
        weight_rom[7484] = 16;
        weight_rom[7485] = 8;
        weight_rom[7486] = 19;
        weight_rom[7487] = 26;
        weight_rom[7488] = 5;
        weight_rom[7489] = -12;
        weight_rom[7490] = -8;
        weight_rom[7491] = 37;
        weight_rom[7492] = 52;
        weight_rom[7493] = 59;
        weight_rom[7494] = 44;
        weight_rom[7495] = 47;
        weight_rom[7496] = 24;
        weight_rom[7497] = 26;
        weight_rom[7498] = 18;
        weight_rom[7499] = -19;
        weight_rom[7500] = 1;
        weight_rom[7501] = 9;
        weight_rom[7502] = 45;
        weight_rom[7503] = 13;
        weight_rom[7504] = -1;
        weight_rom[7505] = 4;
        weight_rom[7506] = -20;
        weight_rom[7507] = -4;
        weight_rom[7508] = 0;
        weight_rom[7509] = 16;
        weight_rom[7510] = 29;
        weight_rom[7511] = 31;
        weight_rom[7512] = 24;
        weight_rom[7513] = 10;
        weight_rom[7514] = 26;
        weight_rom[7515] = 21;
        weight_rom[7516] = 7;
        weight_rom[7517] = -8;
        weight_rom[7518] = 9;
        weight_rom[7519] = 48;
        weight_rom[7520] = 53;
        weight_rom[7521] = 62;
        weight_rom[7522] = 49;
        weight_rom[7523] = 36;
        weight_rom[7524] = 26;
        weight_rom[7525] = 22;
        weight_rom[7526] = 12;
        weight_rom[7527] = -15;
        weight_rom[7528] = 4;
        weight_rom[7529] = 57;
        weight_rom[7530] = 36;
        weight_rom[7531] = 13;
        weight_rom[7532] = 1;
        weight_rom[7533] = -1;
        weight_rom[7534] = 22;
        weight_rom[7535] = -9;
        weight_rom[7536] = -5;
        weight_rom[7537] = 0;
        weight_rom[7538] = 22;
        weight_rom[7539] = 16;
        weight_rom[7540] = 21;
        weight_rom[7541] = 0;
        weight_rom[7542] = 14;
        weight_rom[7543] = 5;
        weight_rom[7544] = 2;
        weight_rom[7545] = 15;
        weight_rom[7546] = 27;
        weight_rom[7547] = 53;
        weight_rom[7548] = 40;
        weight_rom[7549] = 37;
        weight_rom[7550] = 40;
        weight_rom[7551] = 21;
        weight_rom[7552] = 27;
        weight_rom[7553] = 11;
        weight_rom[7554] = 2;
        weight_rom[7555] = -5;
        weight_rom[7556] = 8;
        weight_rom[7557] = 54;
        weight_rom[7558] = 27;
        weight_rom[7559] = 4;
        weight_rom[7560] = -2;
        weight_rom[7561] = 2;
        weight_rom[7562] = -13;
        weight_rom[7563] = -11;
        weight_rom[7564] = 4;
        weight_rom[7565] = -1;
        weight_rom[7566] = 8;
        weight_rom[7567] = 15;
        weight_rom[7568] = 1;
        weight_rom[7569] = -16;
        weight_rom[7570] = -17;
        weight_rom[7571] = -11;
        weight_rom[7572] = -7;
        weight_rom[7573] = 15;
        weight_rom[7574] = 33;
        weight_rom[7575] = 29;
        weight_rom[7576] = 29;
        weight_rom[7577] = 27;
        weight_rom[7578] = 19;
        weight_rom[7579] = 11;
        weight_rom[7580] = 11;
        weight_rom[7581] = 3;
        weight_rom[7582] = -24;
        weight_rom[7583] = -6;
        weight_rom[7584] = 16;
        weight_rom[7585] = 56;
        weight_rom[7586] = 24;
        weight_rom[7587] = 12;
        weight_rom[7588] = 0;
        weight_rom[7589] = 4;
        weight_rom[7590] = 6;
        weight_rom[7591] = 13;
        weight_rom[7592] = 19;
        weight_rom[7593] = -11;
        weight_rom[7594] = -19;
        weight_rom[7595] = -3;
        weight_rom[7596] = -17;
        weight_rom[7597] = -35;
        weight_rom[7598] = -33;
        weight_rom[7599] = -9;
        weight_rom[7600] = 1;
        weight_rom[7601] = 10;
        weight_rom[7602] = 21;
        weight_rom[7603] = 11;
        weight_rom[7604] = 11;
        weight_rom[7605] = -3;
        weight_rom[7606] = -15;
        weight_rom[7607] = -9;
        weight_rom[7608] = -10;
        weight_rom[7609] = -10;
        weight_rom[7610] = -15;
        weight_rom[7611] = -13;
        weight_rom[7612] = -16;
        weight_rom[7613] = 16;
        weight_rom[7614] = 32;
        weight_rom[7615] = 1;
        weight_rom[7616] = -4;
        weight_rom[7617] = -17;
        weight_rom[7618] = 8;
        weight_rom[7619] = 18;
        weight_rom[7620] = 14;
        weight_rom[7621] = -17;
        weight_rom[7622] = -28;
        weight_rom[7623] = -13;
        weight_rom[7624] = -34;
        weight_rom[7625] = -32;
        weight_rom[7626] = -38;
        weight_rom[7627] = -16;
        weight_rom[7628] = 5;
        weight_rom[7629] = -2;
        weight_rom[7630] = 14;
        weight_rom[7631] = -3;
        weight_rom[7632] = -8;
        weight_rom[7633] = -28;
        weight_rom[7634] = -27;
        weight_rom[7635] = -29;
        weight_rom[7636] = -33;
        weight_rom[7637] = -36;
        weight_rom[7638] = -31;
        weight_rom[7639] = -25;
        weight_rom[7640] = 20;
        weight_rom[7641] = -6;
        weight_rom[7642] = 20;
        weight_rom[7643] = 2;
        weight_rom[7644] = -2;
        weight_rom[7645] = 8;
        weight_rom[7646] = 3;
        weight_rom[7647] = -13;
        weight_rom[7648] = -13;
        weight_rom[7649] = -27;
        weight_rom[7650] = -42;
        weight_rom[7651] = -43;
        weight_rom[7652] = -24;
        weight_rom[7653] = -13;
        weight_rom[7654] = -12;
        weight_rom[7655] = 2;
        weight_rom[7656] = 12;
        weight_rom[7657] = 0;
        weight_rom[7658] = -3;
        weight_rom[7659] = -27;
        weight_rom[7660] = -19;
        weight_rom[7661] = -34;
        weight_rom[7662] = -49;
        weight_rom[7663] = -50;
        weight_rom[7664] = -37;
        weight_rom[7665] = -26;
        weight_rom[7666] = -30;
        weight_rom[7667] = -14;
        weight_rom[7668] = 16;
        weight_rom[7669] = -17;
        weight_rom[7670] = 6;
        weight_rom[7671] = 0;
        weight_rom[7672] = 0;
        weight_rom[7673] = 1;
        weight_rom[7674] = -16;
        weight_rom[7675] = -13;
        weight_rom[7676] = -7;
        weight_rom[7677] = -36;
        weight_rom[7678] = -35;
        weight_rom[7679] = -31;
        weight_rom[7680] = -11;
        weight_rom[7681] = 0;
        weight_rom[7682] = 0;
        weight_rom[7683] = 2;
        weight_rom[7684] = -1;
        weight_rom[7685] = -12;
        weight_rom[7686] = -18;
        weight_rom[7687] = -25;
        weight_rom[7688] = -27;
        weight_rom[7689] = -43;
        weight_rom[7690] = -53;
        weight_rom[7691] = -47;
        weight_rom[7692] = -42;
        weight_rom[7693] = -21;
        weight_rom[7694] = -17;
        weight_rom[7695] = -6;
        weight_rom[7696] = 3;
        weight_rom[7697] = -12;
        weight_rom[7698] = -1;
        weight_rom[7699] = -1;
        weight_rom[7700] = 3;
        weight_rom[7701] = 0;
        weight_rom[7702] = -15;
        weight_rom[7703] = -31;
        weight_rom[7704] = -41;
        weight_rom[7705] = -26;
        weight_rom[7706] = -11;
        weight_rom[7707] = 3;
        weight_rom[7708] = -4;
        weight_rom[7709] = -16;
        weight_rom[7710] = -11;
        weight_rom[7711] = -7;
        weight_rom[7712] = -21;
        weight_rom[7713] = -23;
        weight_rom[7714] = -17;
        weight_rom[7715] = -27;
        weight_rom[7716] = -36;
        weight_rom[7717] = -34;
        weight_rom[7718] = -30;
        weight_rom[7719] = -33;
        weight_rom[7720] = -18;
        weight_rom[7721] = 5;
        weight_rom[7722] = -4;
        weight_rom[7723] = -6;
        weight_rom[7724] = 3;
        weight_rom[7725] = -3;
        weight_rom[7726] = -3;
        weight_rom[7727] = 3;
        weight_rom[7728] = 0;
        weight_rom[7729] = -3;
        weight_rom[7730] = -9;
        weight_rom[7731] = -22;
        weight_rom[7732] = -26;
        weight_rom[7733] = 11;
        weight_rom[7734] = 15;
        weight_rom[7735] = 19;
        weight_rom[7736] = 10;
        weight_rom[7737] = -3;
        weight_rom[7738] = -6;
        weight_rom[7739] = -20;
        weight_rom[7740] = -20;
        weight_rom[7741] = -18;
        weight_rom[7742] = -21;
        weight_rom[7743] = -11;
        weight_rom[7744] = -13;
        weight_rom[7745] = 2;
        weight_rom[7746] = -11;
        weight_rom[7747] = -21;
        weight_rom[7748] = 9;
        weight_rom[7749] = 11;
        weight_rom[7750] = 5;
        weight_rom[7751] = -7;
        weight_rom[7752] = 6;
        weight_rom[7753] = 20;
        weight_rom[7754] = -1;
        weight_rom[7755] = -4;
        weight_rom[7756] = -1;
        weight_rom[7757] = 3;
        weight_rom[7758] = 4;
        weight_rom[7759] = -6;
        weight_rom[7760] = -18;
        weight_rom[7761] = 14;
        weight_rom[7762] = 0;
        weight_rom[7763] = 11;
        weight_rom[7764] = 1;
        weight_rom[7765] = 10;
        weight_rom[7766] = 8;
        weight_rom[7767] = 12;
        weight_rom[7768] = 9;
        weight_rom[7769] = 13;
        weight_rom[7770] = 12;
        weight_rom[7771] = 11;
        weight_rom[7772] = 6;
        weight_rom[7773] = 0;
        weight_rom[7774] = 0;
        weight_rom[7775] = -11;
        weight_rom[7776] = 10;
        weight_rom[7777] = 8;
        weight_rom[7778] = -17;
        weight_rom[7779] = -20;
        weight_rom[7780] = -15;
        weight_rom[7781] = -4;
        weight_rom[7782] = -4;
        weight_rom[7783] = 0;
        weight_rom[7784] = 1;
        weight_rom[7785] = 4;
        weight_rom[7786] = -2;
        weight_rom[7787] = 0;
        weight_rom[7788] = 19;
        weight_rom[7789] = 31;
        weight_rom[7790] = 21;
        weight_rom[7791] = 21;
        weight_rom[7792] = 32;
        weight_rom[7793] = 20;
        weight_rom[7794] = 27;
        weight_rom[7795] = 13;
        weight_rom[7796] = 11;
        weight_rom[7797] = 11;
        weight_rom[7798] = 29;
        weight_rom[7799] = 16;
        weight_rom[7800] = 16;
        weight_rom[7801] = 9;
        weight_rom[7802] = 9;
        weight_rom[7803] = 6;
        weight_rom[7804] = 9;
        weight_rom[7805] = 17;
        weight_rom[7806] = 7;
        weight_rom[7807] = 21;
        weight_rom[7808] = -1;
        weight_rom[7809] = -4;
        weight_rom[7810] = -2;
        weight_rom[7811] = 0;
        weight_rom[7812] = -1;
        weight_rom[7813] = -2;
        weight_rom[7814] = -2;
        weight_rom[7815] = 1;
        weight_rom[7816] = -2;
        weight_rom[7817] = 13;
        weight_rom[7818] = 3;
        weight_rom[7819] = 8;
        weight_rom[7820] = 6;
        weight_rom[7821] = 20;
        weight_rom[7822] = 23;
        weight_rom[7823] = 0;
        weight_rom[7824] = 13;
        weight_rom[7825] = 30;
        weight_rom[7826] = 41;
        weight_rom[7827] = 37;
        weight_rom[7828] = 41;
        weight_rom[7829] = 34;
        weight_rom[7830] = 30;
        weight_rom[7831] = 16;
        weight_rom[7832] = 13;
        weight_rom[7833] = 13;
        weight_rom[7834] = 27;
        weight_rom[7835] = 3;
        weight_rom[7836] = 3;
        weight_rom[7837] = 0;
        weight_rom[7838] = 4;
        weight_rom[7839] = 2;
        weight_rom[7840] = -1;
        weight_rom[7841] = 4;
        weight_rom[7842] = -5;
        weight_rom[7843] = 2;
        weight_rom[7844] = 4;
        weight_rom[7845] = -3;
        weight_rom[7846] = -3;
        weight_rom[7847] = 2;
        weight_rom[7848] = 1;
        weight_rom[7849] = -4;
        weight_rom[7850] = 0;
        weight_rom[7851] = 3;
        weight_rom[7852] = -3;
        weight_rom[7853] = -3;
        weight_rom[7854] = 3;
        weight_rom[7855] = -4;
        weight_rom[7856] = 0;
        weight_rom[7857] = 4;
        weight_rom[7858] = 3;
        weight_rom[7859] = 3;
        weight_rom[7860] = -4;
        weight_rom[7861] = -4;
        weight_rom[7862] = -1;
        weight_rom[7863] = 4;
        weight_rom[7864] = -4;
        weight_rom[7865] = 4;
        weight_rom[7866] = -1;
        weight_rom[7867] = -1;
        weight_rom[7868] = -2;
        weight_rom[7869] = 0;
        weight_rom[7870] = 3;
        weight_rom[7871] = 3;
        weight_rom[7872] = 0;
        weight_rom[7873] = -1;
        weight_rom[7874] = 0;
        weight_rom[7875] = -8;
        weight_rom[7876] = -3;
        weight_rom[7877] = -23;
        weight_rom[7878] = -22;
        weight_rom[7879] = -26;
        weight_rom[7880] = -30;
        weight_rom[7881] = -20;
        weight_rom[7882] = 9;
        weight_rom[7883] = 20;
        weight_rom[7884] = 18;
        weight_rom[7885] = -3;
        weight_rom[7886] = -16;
        weight_rom[7887] = -5;
        weight_rom[7888] = -16;
        weight_rom[7889] = -1;
        weight_rom[7890] = 2;
        weight_rom[7891] = 4;
        weight_rom[7892] = -1;
        weight_rom[7893] = 0;
        weight_rom[7894] = 4;
        weight_rom[7895] = -1;
        weight_rom[7896] = 2;
        weight_rom[7897] = -1;
        weight_rom[7898] = 0;
        weight_rom[7899] = -4;
        weight_rom[7900] = -16;
        weight_rom[7901] = -1;
        weight_rom[7902] = -8;
        weight_rom[7903] = -8;
        weight_rom[7904] = -7;
        weight_rom[7905] = 21;
        weight_rom[7906] = -6;
        weight_rom[7907] = 0;
        weight_rom[7908] = 1;
        weight_rom[7909] = 16;
        weight_rom[7910] = 17;
        weight_rom[7911] = 37;
        weight_rom[7912] = 30;
        weight_rom[7913] = 18;
        weight_rom[7914] = 3;
        weight_rom[7915] = -7;
        weight_rom[7916] = -6;
        weight_rom[7917] = 4;
        weight_rom[7918] = -5;
        weight_rom[7919] = -5;
        weight_rom[7920] = 8;
        weight_rom[7921] = 14;
        weight_rom[7922] = 4;
        weight_rom[7923] = -2;
        weight_rom[7924] = -2;
        weight_rom[7925] = 1;
        weight_rom[7926] = -6;
        weight_rom[7927] = 0;
        weight_rom[7928] = 2;
        weight_rom[7929] = -18;
        weight_rom[7930] = -6;
        weight_rom[7931] = -9;
        weight_rom[7932] = -6;
        weight_rom[7933] = 18;
        weight_rom[7934] = 0;
        weight_rom[7935] = -21;
        weight_rom[7936] = -11;
        weight_rom[7937] = 6;
        weight_rom[7938] = -13;
        weight_rom[7939] = -12;
        weight_rom[7940] = -1;
        weight_rom[7941] = -7;
        weight_rom[7942] = -6;
        weight_rom[7943] = -7;
        weight_rom[7944] = -11;
        weight_rom[7945] = 10;
        weight_rom[7946] = 17;
        weight_rom[7947] = -10;
        weight_rom[7948] = -4;
        weight_rom[7949] = 23;
        weight_rom[7950] = 3;
        weight_rom[7951] = 1;
        weight_rom[7952] = -4;
        weight_rom[7953] = 0;
        weight_rom[7954] = 8;
        weight_rom[7955] = 0;
        weight_rom[7956] = -16;
        weight_rom[7957] = -16;
        weight_rom[7958] = -7;
        weight_rom[7959] = -18;
        weight_rom[7960] = -7;
        weight_rom[7961] = -3;
        weight_rom[7962] = -7;
        weight_rom[7963] = -9;
        weight_rom[7964] = 0;
        weight_rom[7965] = 8;
        weight_rom[7966] = 11;
        weight_rom[7967] = 2;
        weight_rom[7968] = 5;
        weight_rom[7969] = 6;
        weight_rom[7970] = 6;
        weight_rom[7971] = -3;
        weight_rom[7972] = 6;
        weight_rom[7973] = -2;
        weight_rom[7974] = -5;
        weight_rom[7975] = 7;
        weight_rom[7976] = 12;
        weight_rom[7977] = 16;
        weight_rom[7978] = 6;
        weight_rom[7979] = -2;
        weight_rom[7980] = -2;
        weight_rom[7981] = -4;
        weight_rom[7982] = -3;
        weight_rom[7983] = -11;
        weight_rom[7984] = -23;
        weight_rom[7985] = -17;
        weight_rom[7986] = -22;
        weight_rom[7987] = -26;
        weight_rom[7988] = -26;
        weight_rom[7989] = -20;
        weight_rom[7990] = -19;
        weight_rom[7991] = -7;
        weight_rom[7992] = 0;
        weight_rom[7993] = 3;
        weight_rom[7994] = -1;
        weight_rom[7995] = -2;
        weight_rom[7996] = 4;
        weight_rom[7997] = 11;
        weight_rom[7998] = 11;
        weight_rom[7999] = 13;
        weight_rom[8000] = 19;
        weight_rom[8001] = 22;
        weight_rom[8002] = 15;
        weight_rom[8003] = 21;
        weight_rom[8004] = 18;
        weight_rom[8005] = 14;
        weight_rom[8006] = 13;
        weight_rom[8007] = 0;
        weight_rom[8008] = -1;
        weight_rom[8009] = -1;
        weight_rom[8010] = -12;
        weight_rom[8011] = -24;
        weight_rom[8012] = -29;
        weight_rom[8013] = -28;
        weight_rom[8014] = -47;
        weight_rom[8015] = -33;
        weight_rom[8016] = -35;
        weight_rom[8017] = -18;
        weight_rom[8018] = -27;
        weight_rom[8019] = -13;
        weight_rom[8020] = -3;
        weight_rom[8021] = -2;
        weight_rom[8022] = 1;
        weight_rom[8023] = 3;
        weight_rom[8024] = 8;
        weight_rom[8025] = 4;
        weight_rom[8026] = 9;
        weight_rom[8027] = 5;
        weight_rom[8028] = 5;
        weight_rom[8029] = 3;
        weight_rom[8030] = -2;
        weight_rom[8031] = 3;
        weight_rom[8032] = 40;
        weight_rom[8033] = 39;
        weight_rom[8034] = 23;
        weight_rom[8035] = -5;
        weight_rom[8036] = -1;
        weight_rom[8037] = -15;
        weight_rom[8038] = 6;
        weight_rom[8039] = -33;
        weight_rom[8040] = -31;
        weight_rom[8041] = -55;
        weight_rom[8042] = -48;
        weight_rom[8043] = -38;
        weight_rom[8044] = -24;
        weight_rom[8045] = -26;
        weight_rom[8046] = -8;
        weight_rom[8047] = -12;
        weight_rom[8048] = -3;
        weight_rom[8049] = 6;
        weight_rom[8050] = 8;
        weight_rom[8051] = 5;
        weight_rom[8052] = 11;
        weight_rom[8053] = -3;
        weight_rom[8054] = 0;
        weight_rom[8055] = -1;
        weight_rom[8056] = 6;
        weight_rom[8057] = -1;
        weight_rom[8058] = 7;
        weight_rom[8059] = 0;
        weight_rom[8060] = -4;
        weight_rom[8061] = 28;
        weight_rom[8062] = 13;
        weight_rom[8063] = 8;
        weight_rom[8064] = -6;
        weight_rom[8065] = -5;
        weight_rom[8066] = -4;
        weight_rom[8067] = -30;
        weight_rom[8068] = -58;
        weight_rom[8069] = -48;
        weight_rom[8070] = -41;
        weight_rom[8071] = -31;
        weight_rom[8072] = -18;
        weight_rom[8073] = -28;
        weight_rom[8074] = -10;
        weight_rom[8075] = -3;
        weight_rom[8076] = 1;
        weight_rom[8077] = 19;
        weight_rom[8078] = 12;
        weight_rom[8079] = 4;
        weight_rom[8080] = -3;
        weight_rom[8081] = -9;
        weight_rom[8082] = -15;
        weight_rom[8083] = -7;
        weight_rom[8084] = -13;
        weight_rom[8085] = 0;
        weight_rom[8086] = -7;
        weight_rom[8087] = 8;
        weight_rom[8088] = 16;
        weight_rom[8089] = 30;
        weight_rom[8090] = 32;
        weight_rom[8091] = 10;
        weight_rom[8092] = 4;
        weight_rom[8093] = -4;
        weight_rom[8094] = -24;
        weight_rom[8095] = -21;
        weight_rom[8096] = -44;
        weight_rom[8097] = -37;
        weight_rom[8098] = -17;
        weight_rom[8099] = -19;
        weight_rom[8100] = -11;
        weight_rom[8101] = -8;
        weight_rom[8102] = 0;
        weight_rom[8103] = 16;
        weight_rom[8104] = 19;
        weight_rom[8105] = 15;
        weight_rom[8106] = 6;
        weight_rom[8107] = 9;
        weight_rom[8108] = -3;
        weight_rom[8109] = -16;
        weight_rom[8110] = -19;
        weight_rom[8111] = -22;
        weight_rom[8112] = -15;
        weight_rom[8113] = -8;
        weight_rom[8114] = -4;
        weight_rom[8115] = 2;
        weight_rom[8116] = 30;
        weight_rom[8117] = 43;
        weight_rom[8118] = 13;
        weight_rom[8119] = -17;
        weight_rom[8120] = -7;
        weight_rom[8121] = -8;
        weight_rom[8122] = -17;
        weight_rom[8123] = -16;
        weight_rom[8124] = -23;
        weight_rom[8125] = -8;
        weight_rom[8126] = -2;
        weight_rom[8127] = -12;
        weight_rom[8128] = -7;
        weight_rom[8129] = 3;
        weight_rom[8130] = 11;
        weight_rom[8131] = 22;
        weight_rom[8132] = 30;
        weight_rom[8133] = 12;
        weight_rom[8134] = 7;
        weight_rom[8135] = 11;
        weight_rom[8136] = -17;
        weight_rom[8137] = -25;
        weight_rom[8138] = -27;
        weight_rom[8139] = -25;
        weight_rom[8140] = -23;
        weight_rom[8141] = -7;
        weight_rom[8142] = -10;
        weight_rom[8143] = -5;
        weight_rom[8144] = 15;
        weight_rom[8145] = 48;
        weight_rom[8146] = 33;
        weight_rom[8147] = 10;
        weight_rom[8148] = -12;
        weight_rom[8149] = -17;
        weight_rom[8150] = -23;
        weight_rom[8151] = -26;
        weight_rom[8152] = -15;
        weight_rom[8153] = 20;
        weight_rom[8154] = 3;
        weight_rom[8155] = 4;
        weight_rom[8156] = 9;
        weight_rom[8157] = 1;
        weight_rom[8158] = 4;
        weight_rom[8159] = 14;
        weight_rom[8160] = 6;
        weight_rom[8161] = 11;
        weight_rom[8162] = 7;
        weight_rom[8163] = -5;
        weight_rom[8164] = -8;
        weight_rom[8165] = -24;
        weight_rom[8166] = -14;
        weight_rom[8167] = -13;
        weight_rom[8168] = -21;
        weight_rom[8169] = -10;
        weight_rom[8170] = -26;
        weight_rom[8171] = -15;
        weight_rom[8172] = 9;
        weight_rom[8173] = 35;
        weight_rom[8174] = 39;
        weight_rom[8175] = 5;
        weight_rom[8176] = -4;
        weight_rom[8177] = -8;
        weight_rom[8178] = -23;
        weight_rom[8179] = -15;
        weight_rom[8180] = 25;
        weight_rom[8181] = 23;
        weight_rom[8182] = 15;
        weight_rom[8183] = 1;
        weight_rom[8184] = 11;
        weight_rom[8185] = 3;
        weight_rom[8186] = 3;
        weight_rom[8187] = 0;
        weight_rom[8188] = 3;
        weight_rom[8189] = 13;
        weight_rom[8190] = 15;
        weight_rom[8191] = 5;
        weight_rom[8192] = -10;
        weight_rom[8193] = -21;
        weight_rom[8194] = -16;
        weight_rom[8195] = -6;
        weight_rom[8196] = -1;
        weight_rom[8197] = -12;
        weight_rom[8198] = -28;
        weight_rom[8199] = -44;
        weight_rom[8200] = -38;
        weight_rom[8201] = 13;
        weight_rom[8202] = 30;
        weight_rom[8203] = 3;
        weight_rom[8204] = 1;
        weight_rom[8205] = 4;
        weight_rom[8206] = -22;
        weight_rom[8207] = 3;
        weight_rom[8208] = 1;
        weight_rom[8209] = 4;
        weight_rom[8210] = 4;
        weight_rom[8211] = 6;
        weight_rom[8212] = 22;
        weight_rom[8213] = 6;
        weight_rom[8214] = 1;
        weight_rom[8215] = 1;
        weight_rom[8216] = 16;
        weight_rom[8217] = 23;
        weight_rom[8218] = 29;
        weight_rom[8219] = 17;
        weight_rom[8220] = -2;
        weight_rom[8221] = -13;
        weight_rom[8222] = -9;
        weight_rom[8223] = -7;
        weight_rom[8224] = -7;
        weight_rom[8225] = -15;
        weight_rom[8226] = -28;
        weight_rom[8227] = -53;
        weight_rom[8228] = -51;
        weight_rom[8229] = 0;
        weight_rom[8230] = 41;
        weight_rom[8231] = 26;
        weight_rom[8232] = -3;
        weight_rom[8233] = -1;
        weight_rom[8234] = 0;
        weight_rom[8235] = 8;
        weight_rom[8236] = 21;
        weight_rom[8237] = 7;
        weight_rom[8238] = 21;
        weight_rom[8239] = 13;
        weight_rom[8240] = 16;
        weight_rom[8241] = 9;
        weight_rom[8242] = -8;
        weight_rom[8243] = 3;
        weight_rom[8244] = 7;
        weight_rom[8245] = 25;
        weight_rom[8246] = 30;
        weight_rom[8247] = 19;
        weight_rom[8248] = 18;
        weight_rom[8249] = -13;
        weight_rom[8250] = -11;
        weight_rom[8251] = -23;
        weight_rom[8252] = -24;
        weight_rom[8253] = -32;
        weight_rom[8254] = -41;
        weight_rom[8255] = -50;
        weight_rom[8256] = -35;
        weight_rom[8257] = 14;
        weight_rom[8258] = 43;
        weight_rom[8259] = 4;
        weight_rom[8260] = 3;
        weight_rom[8261] = -5;
        weight_rom[8262] = -10;
        weight_rom[8263] = 29;
        weight_rom[8264] = 16;
        weight_rom[8265] = 7;
        weight_rom[8266] = 32;
        weight_rom[8267] = 15;
        weight_rom[8268] = 15;
        weight_rom[8269] = 14;
        weight_rom[8270] = 3;
        weight_rom[8271] = -1;
        weight_rom[8272] = 12;
        weight_rom[8273] = 37;
        weight_rom[8274] = 34;
        weight_rom[8275] = 18;
        weight_rom[8276] = 11;
        weight_rom[8277] = -10;
        weight_rom[8278] = -17;
        weight_rom[8279] = -29;
        weight_rom[8280] = -47;
        weight_rom[8281] = -44;
        weight_rom[8282] = -46;
        weight_rom[8283] = -49;
        weight_rom[8284] = -13;
        weight_rom[8285] = 35;
        weight_rom[8286] = 52;
        weight_rom[8287] = 13;
        weight_rom[8288] = -3;
        weight_rom[8289] = 2;
        weight_rom[8290] = -25;
        weight_rom[8291] = 22;
        weight_rom[8292] = 18;
        weight_rom[8293] = 16;
        weight_rom[8294] = 20;
        weight_rom[8295] = 5;
        weight_rom[8296] = -3;
        weight_rom[8297] = 2;
        weight_rom[8298] = 10;
        weight_rom[8299] = 16;
        weight_rom[8300] = 29;
        weight_rom[8301] = 33;
        weight_rom[8302] = 34;
        weight_rom[8303] = 17;
        weight_rom[8304] = 10;
        weight_rom[8305] = -8;
        weight_rom[8306] = -31;
        weight_rom[8307] = -39;
        weight_rom[8308] = -34;
        weight_rom[8309] = -27;
        weight_rom[8310] = -14;
        weight_rom[8311] = -21;
        weight_rom[8312] = 3;
        weight_rom[8313] = 62;
        weight_rom[8314] = 61;
        weight_rom[8315] = 25;
        weight_rom[8316] = 4;
        weight_rom[8317] = -8;
        weight_rom[8318] = 10;
        weight_rom[8319] = 9;
        weight_rom[8320] = -4;
        weight_rom[8321] = 15;
        weight_rom[8322] = 18;
        weight_rom[8323] = -3;
        weight_rom[8324] = 2;
        weight_rom[8325] = 8;
        weight_rom[8326] = 23;
        weight_rom[8327] = 23;
        weight_rom[8328] = 25;
        weight_rom[8329] = 29;
        weight_rom[8330] = 23;
        weight_rom[8331] = 22;
        weight_rom[8332] = -5;
        weight_rom[8333] = -20;
        weight_rom[8334] = -25;
        weight_rom[8335] = -29;
        weight_rom[8336] = -10;
        weight_rom[8337] = -16;
        weight_rom[8338] = -16;
        weight_rom[8339] = -20;
        weight_rom[8340] = 6;
        weight_rom[8341] = 40;
        weight_rom[8342] = 59;
        weight_rom[8343] = 3;
        weight_rom[8344] = -4;
        weight_rom[8345] = -6;
        weight_rom[8346] = -6;
        weight_rom[8347] = 3;
        weight_rom[8348] = 1;
        weight_rom[8349] = 12;
        weight_rom[8350] = 10;
        weight_rom[8351] = 7;
        weight_rom[8352] = 6;
        weight_rom[8353] = 14;
        weight_rom[8354] = 19;
        weight_rom[8355] = 24;
        weight_rom[8356] = 23;
        weight_rom[8357] = 24;
        weight_rom[8358] = 32;
        weight_rom[8359] = 3;
        weight_rom[8360] = -6;
        weight_rom[8361] = -10;
        weight_rom[8362] = -12;
        weight_rom[8363] = -4;
        weight_rom[8364] = 4;
        weight_rom[8365] = -1;
        weight_rom[8366] = -7;
        weight_rom[8367] = 8;
        weight_rom[8368] = 40;
        weight_rom[8369] = 56;
        weight_rom[8370] = 27;
        weight_rom[8371] = 22;
        weight_rom[8372] = -4;
        weight_rom[8373] = -1;
        weight_rom[8374] = -3;
        weight_rom[8375] = -23;
        weight_rom[8376] = -1;
        weight_rom[8377] = -10;
        weight_rom[8378] = 2;
        weight_rom[8379] = 3;
        weight_rom[8380] = 6;
        weight_rom[8381] = 21;
        weight_rom[8382] = 10;
        weight_rom[8383] = 11;
        weight_rom[8384] = 2;
        weight_rom[8385] = 22;
        weight_rom[8386] = 7;
        weight_rom[8387] = 6;
        weight_rom[8388] = 6;
        weight_rom[8389] = 1;
        weight_rom[8390] = 10;
        weight_rom[8391] = 10;
        weight_rom[8392] = 12;
        weight_rom[8393] = 5;
        weight_rom[8394] = 6;
        weight_rom[8395] = 16;
        weight_rom[8396] = 21;
        weight_rom[8397] = 54;
        weight_rom[8398] = 37;
        weight_rom[8399] = 12;
        weight_rom[8400] = 4;
        weight_rom[8401] = -18;
        weight_rom[8402] = 10;
        weight_rom[8403] = -5;
        weight_rom[8404] = -7;
        weight_rom[8405] = -4;
        weight_rom[8406] = 1;
        weight_rom[8407] = 1;
        weight_rom[8408] = 7;
        weight_rom[8409] = 9;
        weight_rom[8410] = 4;
        weight_rom[8411] = 1;
        weight_rom[8412] = -6;
        weight_rom[8413] = -12;
        weight_rom[8414] = -5;
        weight_rom[8415] = 5;
        weight_rom[8416] = 17;
        weight_rom[8417] = 20;
        weight_rom[8418] = 30;
        weight_rom[8419] = 21;
        weight_rom[8420] = 22;
        weight_rom[8421] = 22;
        weight_rom[8422] = 30;
        weight_rom[8423] = 30;
        weight_rom[8424] = 48;
        weight_rom[8425] = 48;
        weight_rom[8426] = 21;
        weight_rom[8427] = -2;
        weight_rom[8428] = -3;
        weight_rom[8429] = 13;
        weight_rom[8430] = -18;
        weight_rom[8431] = -4;
        weight_rom[8432] = 8;
        weight_rom[8433] = 6;
        weight_rom[8434] = -1;
        weight_rom[8435] = -5;
        weight_rom[8436] = -3;
        weight_rom[8437] = 5;
        weight_rom[8438] = -6;
        weight_rom[8439] = -9;
        weight_rom[8440] = -11;
        weight_rom[8441] = -8;
        weight_rom[8442] = -6;
        weight_rom[8443] = 2;
        weight_rom[8444] = 4;
        weight_rom[8445] = 22;
        weight_rom[8446] = 22;
        weight_rom[8447] = 29;
        weight_rom[8448] = 32;
        weight_rom[8449] = 34;
        weight_rom[8450] = 42;
        weight_rom[8451] = 59;
        weight_rom[8452] = 61;
        weight_rom[8453] = 40;
        weight_rom[8454] = -3;
        weight_rom[8455] = -4;
        weight_rom[8456] = -1;
        weight_rom[8457] = 4;
        weight_rom[8458] = -15;
        weight_rom[8459] = 6;
        weight_rom[8460] = 24;
        weight_rom[8461] = 17;
        weight_rom[8462] = 0;
        weight_rom[8463] = -3;
        weight_rom[8464] = -2;
        weight_rom[8465] = -7;
        weight_rom[8466] = -3;
        weight_rom[8467] = -6;
        weight_rom[8468] = -16;
        weight_rom[8469] = -17;
        weight_rom[8470] = 2;
        weight_rom[8471] = -1;
        weight_rom[8472] = -4;
        weight_rom[8473] = 15;
        weight_rom[8474] = 31;
        weight_rom[8475] = 22;
        weight_rom[8476] = 41;
        weight_rom[8477] = 30;
        weight_rom[8478] = 38;
        weight_rom[8479] = 36;
        weight_rom[8480] = 56;
        weight_rom[8481] = 31;
        weight_rom[8482] = 6;
        weight_rom[8483] = -3;
        weight_rom[8484] = 0;
        weight_rom[8485] = 0;
        weight_rom[8486] = -1;
        weight_rom[8487] = -17;
        weight_rom[8488] = -5;
        weight_rom[8489] = -9;
        weight_rom[8490] = -23;
        weight_rom[8491] = -27;
        weight_rom[8492] = -8;
        weight_rom[8493] = -9;
        weight_rom[8494] = -14;
        weight_rom[8495] = -8;
        weight_rom[8496] = -3;
        weight_rom[8497] = -2;
        weight_rom[8498] = -6;
        weight_rom[8499] = -4;
        weight_rom[8500] = 10;
        weight_rom[8501] = 7;
        weight_rom[8502] = 16;
        weight_rom[8503] = 27;
        weight_rom[8504] = 37;
        weight_rom[8505] = 30;
        weight_rom[8506] = 51;
        weight_rom[8507] = 38;
        weight_rom[8508] = 39;
        weight_rom[8509] = 19;
        weight_rom[8510] = 9;
        weight_rom[8511] = -3;
        weight_rom[8512] = 1;
        weight_rom[8513] = 1;
        weight_rom[8514] = -4;
        weight_rom[8515] = -39;
        weight_rom[8516] = -22;
        weight_rom[8517] = -46;
        weight_rom[8518] = -35;
        weight_rom[8519] = -39;
        weight_rom[8520] = -20;
        weight_rom[8521] = -6;
        weight_rom[8522] = -20;
        weight_rom[8523] = -17;
        weight_rom[8524] = -12;
        weight_rom[8525] = -10;
        weight_rom[8526] = -3;
        weight_rom[8527] = 3;
        weight_rom[8528] = 1;
        weight_rom[8529] = 17;
        weight_rom[8530] = 38;
        weight_rom[8531] = 37;
        weight_rom[8532] = 30;
        weight_rom[8533] = 32;
        weight_rom[8534] = 34;
        weight_rom[8535] = 27;
        weight_rom[8536] = 25;
        weight_rom[8537] = 15;
        weight_rom[8538] = 4;
        weight_rom[8539] = -2;
        weight_rom[8540] = -1;
        weight_rom[8541] = -1;
        weight_rom[8542] = 2;
        weight_rom[8543] = -8;
        weight_rom[8544] = -23;
        weight_rom[8545] = -35;
        weight_rom[8546] = -34;
        weight_rom[8547] = -17;
        weight_rom[8548] = -20;
        weight_rom[8549] = -20;
        weight_rom[8550] = -17;
        weight_rom[8551] = -13;
        weight_rom[8552] = -6;
        weight_rom[8553] = 7;
        weight_rom[8554] = 13;
        weight_rom[8555] = 3;
        weight_rom[8556] = 18;
        weight_rom[8557] = 22;
        weight_rom[8558] = 5;
        weight_rom[8559] = -1;
        weight_rom[8560] = 17;
        weight_rom[8561] = 18;
        weight_rom[8562] = 6;
        weight_rom[8563] = 37;
        weight_rom[8564] = 33;
        weight_rom[8565] = 2;
        weight_rom[8566] = 0;
        weight_rom[8567] = -4;
        weight_rom[8568] = 1;
        weight_rom[8569] = 3;
        weight_rom[8570] = 3;
        weight_rom[8571] = -2;
        weight_rom[8572] = 17;
        weight_rom[8573] = 9;
        weight_rom[8574] = 1;
        weight_rom[8575] = -2;
        weight_rom[8576] = 11;
        weight_rom[8577] = 1;
        weight_rom[8578] = 7;
        weight_rom[8579] = 28;
        weight_rom[8580] = 38;
        weight_rom[8581] = 14;
        weight_rom[8582] = 22;
        weight_rom[8583] = 16;
        weight_rom[8584] = 6;
        weight_rom[8585] = -2;
        weight_rom[8586] = 7;
        weight_rom[8587] = -16;
        weight_rom[8588] = 1;
        weight_rom[8589] = 4;
        weight_rom[8590] = -3;
        weight_rom[8591] = 5;
        weight_rom[8592] = -1;
        weight_rom[8593] = 2;
        weight_rom[8594] = -1;
        weight_rom[8595] = 4;
        weight_rom[8596] = 2;
        weight_rom[8597] = -3;
        weight_rom[8598] = -2;
        weight_rom[8599] = 1;
        weight_rom[8600] = 3;
        weight_rom[8601] = -1;
        weight_rom[8602] = -9;
        weight_rom[8603] = 10;
        weight_rom[8604] = 7;
        weight_rom[8605] = 6;
        weight_rom[8606] = -3;
        weight_rom[8607] = 24;
        weight_rom[8608] = 20;
        weight_rom[8609] = -21;
        weight_rom[8610] = 15;
        weight_rom[8611] = 21;
        weight_rom[8612] = 5;
        weight_rom[8613] = -40;
        weight_rom[8614] = -20;
        weight_rom[8615] = 5;
        weight_rom[8616] = -5;
        weight_rom[8617] = -7;
        weight_rom[8618] = 3;
        weight_rom[8619] = -4;
        weight_rom[8620] = 0;
        weight_rom[8621] = 2;
        weight_rom[8622] = -4;
        weight_rom[8623] = -4;
        weight_rom[8624] = 1;
        weight_rom[8625] = 3;
        weight_rom[8626] = 3;
        weight_rom[8627] = -2;
        weight_rom[8628] = 3;
        weight_rom[8629] = 0;
        weight_rom[8630] = 3;
        weight_rom[8631] = 3;
        weight_rom[8632] = 1;
        weight_rom[8633] = 2;
        weight_rom[8634] = -2;
        weight_rom[8635] = -2;
        weight_rom[8636] = -4;
        weight_rom[8637] = 6;
        weight_rom[8638] = 3;
        weight_rom[8639] = -4;
        weight_rom[8640] = -2;
        weight_rom[8641] = -4;
        weight_rom[8642] = 4;
        weight_rom[8643] = 2;
        weight_rom[8644] = 0;
        weight_rom[8645] = 0;
        weight_rom[8646] = 1;
        weight_rom[8647] = -2;
        weight_rom[8648] = -2;
        weight_rom[8649] = -1;
        weight_rom[8650] = 4;
        weight_rom[8651] = -1;
        weight_rom[8652] = 4;
        weight_rom[8653] = -2;
        weight_rom[8654] = 0;
        weight_rom[8655] = -2;
        weight_rom[8656] = -1;
        weight_rom[8657] = -1;
        weight_rom[8658] = 11;
        weight_rom[8659] = 13;
        weight_rom[8660] = 25;
        weight_rom[8661] = 8;
        weight_rom[8662] = 11;
        weight_rom[8663] = 13;
        weight_rom[8664] = 25;
        weight_rom[8665] = 26;
        weight_rom[8666] = 4;
        weight_rom[8667] = 1;
        weight_rom[8668] = 33;
        weight_rom[8669] = 16;
        weight_rom[8670] = 20;
        weight_rom[8671] = 21;
        weight_rom[8672] = 11;
        weight_rom[8673] = 9;
        weight_rom[8674] = 7;
        weight_rom[8675] = 4;
        weight_rom[8676] = 4;
        weight_rom[8677] = 3;
        weight_rom[8678] = -1;
        weight_rom[8679] = -5;
        weight_rom[8680] = 4;
        weight_rom[8681] = -3;
        weight_rom[8682] = 2;
        weight_rom[8683] = 0;
        weight_rom[8684] = -3;
        weight_rom[8685] = 3;
        weight_rom[8686] = 8;
        weight_rom[8687] = 18;
        weight_rom[8688] = 30;
        weight_rom[8689] = 36;
        weight_rom[8690] = 41;
        weight_rom[8691] = 35;
        weight_rom[8692] = 28;
        weight_rom[8693] = 11;
        weight_rom[8694] = 11;
        weight_rom[8695] = -10;
        weight_rom[8696] = 21;
        weight_rom[8697] = 35;
        weight_rom[8698] = 59;
        weight_rom[8699] = 18;
        weight_rom[8700] = 20;
        weight_rom[8701] = 20;
        weight_rom[8702] = 9;
        weight_rom[8703] = 15;
        weight_rom[8704] = 11;
        weight_rom[8705] = -4;
        weight_rom[8706] = 1;
        weight_rom[8707] = -1;
        weight_rom[8708] = 2;
        weight_rom[8709] = -1;
        weight_rom[8710] = 8;
        weight_rom[8711] = -3;
        weight_rom[8712] = 0;
        weight_rom[8713] = -4;
        weight_rom[8714] = 7;
        weight_rom[8715] = 1;
        weight_rom[8716] = 25;
        weight_rom[8717] = 34;
        weight_rom[8718] = 37;
        weight_rom[8719] = 46;
        weight_rom[8720] = 47;
        weight_rom[8721] = 33;
        weight_rom[8722] = 15;
        weight_rom[8723] = 10;
        weight_rom[8724] = 5;
        weight_rom[8725] = 32;
        weight_rom[8726] = 37;
        weight_rom[8727] = 30;
        weight_rom[8728] = 41;
        weight_rom[8729] = 42;
        weight_rom[8730] = 36;
        weight_rom[8731] = 27;
        weight_rom[8732] = 28;
        weight_rom[8733] = 15;
        weight_rom[8734] = 4;
        weight_rom[8735] = -2;
        weight_rom[8736] = 2;
        weight_rom[8737] = -2;
        weight_rom[8738] = -11;
        weight_rom[8739] = 0;
        weight_rom[8740] = -1;
        weight_rom[8741] = -14;
        weight_rom[8742] = -27;
        weight_rom[8743] = -8;
        weight_rom[8744] = 2;
        weight_rom[8745] = 32;
        weight_rom[8746] = 44;
        weight_rom[8747] = 38;
        weight_rom[8748] = 28;
        weight_rom[8749] = 12;
        weight_rom[8750] = 22;
        weight_rom[8751] = 22;
        weight_rom[8752] = 13;
        weight_rom[8753] = 22;
        weight_rom[8754] = 30;
        weight_rom[8755] = 15;
        weight_rom[8756] = 5;
        weight_rom[8757] = 20;
        weight_rom[8758] = 0;
        weight_rom[8759] = 7;
        weight_rom[8760] = 15;
        weight_rom[8761] = 8;
        weight_rom[8762] = 14;
        weight_rom[8763] = 1;
        weight_rom[8764] = -1;
        weight_rom[8765] = 1;
        weight_rom[8766] = 3;
        weight_rom[8767] = 0;
        weight_rom[8768] = -11;
        weight_rom[8769] = -31;
        weight_rom[8770] = -17;
        weight_rom[8771] = 0;
        weight_rom[8772] = 1;
        weight_rom[8773] = 18;
        weight_rom[8774] = 32;
        weight_rom[8775] = 28;
        weight_rom[8776] = 13;
        weight_rom[8777] = 14;
        weight_rom[8778] = 10;
        weight_rom[8779] = 11;
        weight_rom[8780] = 20;
        weight_rom[8781] = 21;
        weight_rom[8782] = 21;
        weight_rom[8783] = 14;
        weight_rom[8784] = 28;
        weight_rom[8785] = 20;
        weight_rom[8786] = 13;
        weight_rom[8787] = 4;
        weight_rom[8788] = 7;
        weight_rom[8789] = 29;
        weight_rom[8790] = 14;
        weight_rom[8791] = -1;
        weight_rom[8792] = -1;
        weight_rom[8793] = 4;
        weight_rom[8794] = 2;
        weight_rom[8795] = 11;
        weight_rom[8796] = -1;
        weight_rom[8797] = -1;
        weight_rom[8798] = 3;
        weight_rom[8799] = 10;
        weight_rom[8800] = 12;
        weight_rom[8801] = 14;
        weight_rom[8802] = 11;
        weight_rom[8803] = 7;
        weight_rom[8804] = 13;
        weight_rom[8805] = 21;
        weight_rom[8806] = 18;
        weight_rom[8807] = 23;
        weight_rom[8808] = 22;
        weight_rom[8809] = 19;
        weight_rom[8810] = 15;
        weight_rom[8811] = 10;
        weight_rom[8812] = 11;
        weight_rom[8813] = 12;
        weight_rom[8814] = 17;
        weight_rom[8815] = 7;
        weight_rom[8816] = 39;
        weight_rom[8817] = 39;
        weight_rom[8818] = 12;
        weight_rom[8819] = 11;
        weight_rom[8820] = -1;
        weight_rom[8821] = 13;
        weight_rom[8822] = -17;
        weight_rom[8823] = 0;
        weight_rom[8824] = 9;
        weight_rom[8825] = 5;
        weight_rom[8826] = 5;
        weight_rom[8827] = 5;
        weight_rom[8828] = 25;
        weight_rom[8829] = 10;
        weight_rom[8830] = 11;
        weight_rom[8831] = 13;
        weight_rom[8832] = 13;
        weight_rom[8833] = 15;
        weight_rom[8834] = 18;
        weight_rom[8835] = 23;
        weight_rom[8836] = 21;
        weight_rom[8837] = 10;
        weight_rom[8838] = 10;
        weight_rom[8839] = 7;
        weight_rom[8840] = 9;
        weight_rom[8841] = 4;
        weight_rom[8842] = 10;
        weight_rom[8843] = 7;
        weight_rom[8844] = 16;
        weight_rom[8845] = 15;
        weight_rom[8846] = -4;
        weight_rom[8847] = 6;
        weight_rom[8848] = -9;
        weight_rom[8849] = 4;
        weight_rom[8850] = -10;
        weight_rom[8851] = 6;
        weight_rom[8852] = 1;
        weight_rom[8853] = -3;
        weight_rom[8854] = 8;
        weight_rom[8855] = 14;
        weight_rom[8856] = 3;
        weight_rom[8857] = 14;
        weight_rom[8858] = 22;
        weight_rom[8859] = 11;
        weight_rom[8860] = 23;
        weight_rom[8861] = 19;
        weight_rom[8862] = 25;
        weight_rom[8863] = 8;
        weight_rom[8864] = 19;
        weight_rom[8865] = 7;
        weight_rom[8866] = -2;
        weight_rom[8867] = 9;
        weight_rom[8868] = 13;
        weight_rom[8869] = 7;
        weight_rom[8870] = 7;
        weight_rom[8871] = 10;
        weight_rom[8872] = 22;
        weight_rom[8873] = 9;
        weight_rom[8874] = 20;
        weight_rom[8875] = 8;
        weight_rom[8876] = -2;
        weight_rom[8877] = 2;
        weight_rom[8878] = -17;
        weight_rom[8879] = -3;
        weight_rom[8880] = 10;
        weight_rom[8881] = 10;
        weight_rom[8882] = 3;
        weight_rom[8883] = 5;
        weight_rom[8884] = 17;
        weight_rom[8885] = 18;
        weight_rom[8886] = 10;
        weight_rom[8887] = 15;
        weight_rom[8888] = 7;
        weight_rom[8889] = 15;
        weight_rom[8890] = 17;
        weight_rom[8891] = -6;
        weight_rom[8892] = -7;
        weight_rom[8893] = -17;
        weight_rom[8894] = -7;
        weight_rom[8895] = -10;
        weight_rom[8896] = -1;
        weight_rom[8897] = -3;
        weight_rom[8898] = -6;
        weight_rom[8899] = 6;
        weight_rom[8900] = 35;
        weight_rom[8901] = 41;
        weight_rom[8902] = 14;
        weight_rom[8903] = -16;
        weight_rom[8904] = -11;
        weight_rom[8905] = -13;
        weight_rom[8906] = 2;
        weight_rom[8907] = 13;
        weight_rom[8908] = 20;
        weight_rom[8909] = 9;
        weight_rom[8910] = 20;
        weight_rom[8911] = 6;
        weight_rom[8912] = 1;
        weight_rom[8913] = 15;
        weight_rom[8914] = 7;
        weight_rom[8915] = 5;
        weight_rom[8916] = 5;
        weight_rom[8917] = 17;
        weight_rom[8918] = 8;
        weight_rom[8919] = -21;
        weight_rom[8920] = -26;
        weight_rom[8921] = -28;
        weight_rom[8922] = -21;
        weight_rom[8923] = -26;
        weight_rom[8924] = -13;
        weight_rom[8925] = -20;
        weight_rom[8926] = -20;
        weight_rom[8927] = 9;
        weight_rom[8928] = 41;
        weight_rom[8929] = 32;
        weight_rom[8930] = 19;
        weight_rom[8931] = 10;
        weight_rom[8932] = -19;
        weight_rom[8933] = 0;
        weight_rom[8934] = -8;
        weight_rom[8935] = -6;
        weight_rom[8936] = 20;
        weight_rom[8937] = 9;
        weight_rom[8938] = 12;
        weight_rom[8939] = -1;
        weight_rom[8940] = 3;
        weight_rom[8941] = 2;
        weight_rom[8942] = -9;
        weight_rom[8943] = -5;
        weight_rom[8944] = 2;
        weight_rom[8945] = 23;
        weight_rom[8946] = 16;
        weight_rom[8947] = -37;
        weight_rom[8948] = -42;
        weight_rom[8949] = -29;
        weight_rom[8950] = -21;
        weight_rom[8951] = -28;
        weight_rom[8952] = -42;
        weight_rom[8953] = -44;
        weight_rom[8954] = -42;
        weight_rom[8955] = -15;
        weight_rom[8956] = 21;
        weight_rom[8957] = 26;
        weight_rom[8958] = 35;
        weight_rom[8959] = -14;
        weight_rom[8960] = -11;
        weight_rom[8961] = 0;
        weight_rom[8962] = 5;
        weight_rom[8963] = 7;
        weight_rom[8964] = -4;
        weight_rom[8965] = -12;
        weight_rom[8966] = -8;
        weight_rom[8967] = 0;
        weight_rom[8968] = -4;
        weight_rom[8969] = 0;
        weight_rom[8970] = -6;
        weight_rom[8971] = -5;
        weight_rom[8972] = 3;
        weight_rom[8973] = 15;
        weight_rom[8974] = -9;
        weight_rom[8975] = -19;
        weight_rom[8976] = -33;
        weight_rom[8977] = -21;
        weight_rom[8978] = -20;
        weight_rom[8979] = -24;
        weight_rom[8980] = -19;
        weight_rom[8981] = -38;
        weight_rom[8982] = -53;
        weight_rom[8983] = -39;
        weight_rom[8984] = -7;
        weight_rom[8985] = 30;
        weight_rom[8986] = 32;
        weight_rom[8987] = -8;
        weight_rom[8988] = -4;
        weight_rom[8989] = 2;
        weight_rom[8990] = 7;
        weight_rom[8991] = 10;
        weight_rom[8992] = -34;
        weight_rom[8993] = -21;
        weight_rom[8994] = -11;
        weight_rom[8995] = -15;
        weight_rom[8996] = -8;
        weight_rom[8997] = -5;
        weight_rom[8998] = -13;
        weight_rom[8999] = -5;
        weight_rom[9000] = 10;
        weight_rom[9001] = 11;
        weight_rom[9002] = -7;
        weight_rom[9003] = -17;
        weight_rom[9004] = -23;
        weight_rom[9005] = -22;
        weight_rom[9006] = -15;
        weight_rom[9007] = -4;
        weight_rom[9008] = -21;
        weight_rom[9009] = -34;
        weight_rom[9010] = -27;
        weight_rom[9011] = -26;
        weight_rom[9012] = -8;
        weight_rom[9013] = 8;
        weight_rom[9014] = 20;
        weight_rom[9015] = 17;
        weight_rom[9016] = 1;
        weight_rom[9017] = 1;
        weight_rom[9018] = -8;
        weight_rom[9019] = 1;
        weight_rom[9020] = -26;
        weight_rom[9021] = -31;
        weight_rom[9022] = -18;
        weight_rom[9023] = -8;
        weight_rom[9024] = -8;
        weight_rom[9025] = -12;
        weight_rom[9026] = 3;
        weight_rom[9027] = -1;
        weight_rom[9028] = 9;
        weight_rom[9029] = 10;
        weight_rom[9030] = -5;
        weight_rom[9031] = -12;
        weight_rom[9032] = -22;
        weight_rom[9033] = -16;
        weight_rom[9034] = -18;
        weight_rom[9035] = -24;
        weight_rom[9036] = -15;
        weight_rom[9037] = -18;
        weight_rom[9038] = -27;
        weight_rom[9039] = -14;
        weight_rom[9040] = 10;
        weight_rom[9041] = -3;
        weight_rom[9042] = 12;
        weight_rom[9043] = 0;
        weight_rom[9044] = 2;
        weight_rom[9045] = 0;
        weight_rom[9046] = 8;
        weight_rom[9047] = -8;
        weight_rom[9048] = -19;
        weight_rom[9049] = -23;
        weight_rom[9050] = -15;
        weight_rom[9051] = -15;
        weight_rom[9052] = -11;
        weight_rom[9053] = 1;
        weight_rom[9054] = 7;
        weight_rom[9055] = 1;
        weight_rom[9056] = 10;
        weight_rom[9057] = 12;
        weight_rom[9058] = -4;
        weight_rom[9059] = -14;
        weight_rom[9060] = -19;
        weight_rom[9061] = -15;
        weight_rom[9062] = -10;
        weight_rom[9063] = -9;
        weight_rom[9064] = -9;
        weight_rom[9065] = -20;
        weight_rom[9066] = -23;
        weight_rom[9067] = 2;
        weight_rom[9068] = 33;
        weight_rom[9069] = 20;
        weight_rom[9070] = 1;
        weight_rom[9071] = 3;
        weight_rom[9072] = 1;
        weight_rom[9073] = -2;
        weight_rom[9074] = 3;
        weight_rom[9075] = 13;
        weight_rom[9076] = -22;
        weight_rom[9077] = -35;
        weight_rom[9078] = -38;
        weight_rom[9079] = -40;
        weight_rom[9080] = -17;
        weight_rom[9081] = -2;
        weight_rom[9082] = 6;
        weight_rom[9083] = 18;
        weight_rom[9084] = 20;
        weight_rom[9085] = 11;
        weight_rom[9086] = -2;
        weight_rom[9087] = -16;
        weight_rom[9088] = -18;
        weight_rom[9089] = -11;
        weight_rom[9090] = -13;
        weight_rom[9091] = 5;
        weight_rom[9092] = -6;
        weight_rom[9093] = 7;
        weight_rom[9094] = 19;
        weight_rom[9095] = 20;
        weight_rom[9096] = 38;
        weight_rom[9097] = 28;
        weight_rom[9098] = 13;
        weight_rom[9099] = -6;
        weight_rom[9100] = 0;
        weight_rom[9101] = -9;
        weight_rom[9102] = 3;
        weight_rom[9103] = 13;
        weight_rom[9104] = -15;
        weight_rom[9105] = -23;
        weight_rom[9106] = -30;
        weight_rom[9107] = -47;
        weight_rom[9108] = -38;
        weight_rom[9109] = -16;
        weight_rom[9110] = 5;
        weight_rom[9111] = 9;
        weight_rom[9112] = -1;
        weight_rom[9113] = -15;
        weight_rom[9114] = -31;
        weight_rom[9115] = -23;
        weight_rom[9116] = -13;
        weight_rom[9117] = 3;
        weight_rom[9118] = 7;
        weight_rom[9119] = 11;
        weight_rom[9120] = 7;
        weight_rom[9121] = 12;
        weight_rom[9122] = 22;
        weight_rom[9123] = 25;
        weight_rom[9124] = 21;
        weight_rom[9125] = -1;
        weight_rom[9126] = 9;
        weight_rom[9127] = 4;
        weight_rom[9128] = 3;
        weight_rom[9129] = -4;
        weight_rom[9130] = 17;
        weight_rom[9131] = 10;
        weight_rom[9132] = 1;
        weight_rom[9133] = -3;
        weight_rom[9134] = -21;
        weight_rom[9135] = -39;
        weight_rom[9136] = -34;
        weight_rom[9137] = -26;
        weight_rom[9138] = -11;
        weight_rom[9139] = -9;
        weight_rom[9140] = -9;
        weight_rom[9141] = -23;
        weight_rom[9142] = -32;
        weight_rom[9143] = -20;
        weight_rom[9144] = -2;
        weight_rom[9145] = 10;
        weight_rom[9146] = 2;
        weight_rom[9147] = 18;
        weight_rom[9148] = 4;
        weight_rom[9149] = 8;
        weight_rom[9150] = 32;
        weight_rom[9151] = 22;
        weight_rom[9152] = 27;
        weight_rom[9153] = 6;
        weight_rom[9154] = -9;
        weight_rom[9155] = 1;
        weight_rom[9156] = 1;
        weight_rom[9157] = -11;
        weight_rom[9158] = 11;
        weight_rom[9159] = -2;
        weight_rom[9160] = 22;
        weight_rom[9161] = 10;
        weight_rom[9162] = 6;
        weight_rom[9163] = -6;
        weight_rom[9164] = -1;
        weight_rom[9165] = -8;
        weight_rom[9166] = 7;
        weight_rom[9167] = -14;
        weight_rom[9168] = 1;
        weight_rom[9169] = -5;
        weight_rom[9170] = -10;
        weight_rom[9171] = 2;
        weight_rom[9172] = -1;
        weight_rom[9173] = 16;
        weight_rom[9174] = 16;
        weight_rom[9175] = 14;
        weight_rom[9176] = 22;
        weight_rom[9177] = 23;
        weight_rom[9178] = 31;
        weight_rom[9179] = 27;
        weight_rom[9180] = 2;
        weight_rom[9181] = 3;
        weight_rom[9182] = -10;
        weight_rom[9183] = -8;
        weight_rom[9184] = -3;
        weight_rom[9185] = 9;
        weight_rom[9186] = 6;
        weight_rom[9187] = 16;
        weight_rom[9188] = 7;
        weight_rom[9189] = 31;
        weight_rom[9190] = 15;
        weight_rom[9191] = 18;
        weight_rom[9192] = 21;
        weight_rom[9193] = 17;
        weight_rom[9194] = 19;
        weight_rom[9195] = 1;
        weight_rom[9196] = 15;
        weight_rom[9197] = 16;
        weight_rom[9198] = 5;
        weight_rom[9199] = 10;
        weight_rom[9200] = 9;
        weight_rom[9201] = 10;
        weight_rom[9202] = 19;
        weight_rom[9203] = 6;
        weight_rom[9204] = 20;
        weight_rom[9205] = 35;
        weight_rom[9206] = 38;
        weight_rom[9207] = 31;
        weight_rom[9208] = -8;
        weight_rom[9209] = 7;
        weight_rom[9210] = -14;
        weight_rom[9211] = -2;
        weight_rom[9212] = 0;
        weight_rom[9213] = -9;
        weight_rom[9214] = 18;
        weight_rom[9215] = 23;
        weight_rom[9216] = 16;
        weight_rom[9217] = 15;
        weight_rom[9218] = 22;
        weight_rom[9219] = 24;
        weight_rom[9220] = 22;
        weight_rom[9221] = 15;
        weight_rom[9222] = 8;
        weight_rom[9223] = 23;
        weight_rom[9224] = 30;
        weight_rom[9225] = 30;
        weight_rom[9226] = 28;
        weight_rom[9227] = 27;
        weight_rom[9228] = 15;
        weight_rom[9229] = 12;
        weight_rom[9230] = 10;
        weight_rom[9231] = 12;
        weight_rom[9232] = 7;
        weight_rom[9233] = 12;
        weight_rom[9234] = 42;
        weight_rom[9235] = 37;
        weight_rom[9236] = -6;
        weight_rom[9237] = 9;
        weight_rom[9238] = -7;
        weight_rom[9239] = -1;
        weight_rom[9240] = -1;
        weight_rom[9241] = 4;
        weight_rom[9242] = 21;
        weight_rom[9243] = 20;
        weight_rom[9244] = 6;
        weight_rom[9245] = -5;
        weight_rom[9246] = 13;
        weight_rom[9247] = 29;
        weight_rom[9248] = 22;
        weight_rom[9249] = 17;
        weight_rom[9250] = 13;
        weight_rom[9251] = 22;
        weight_rom[9252] = 32;
        weight_rom[9253] = 30;
        weight_rom[9254] = 23;
        weight_rom[9255] = 24;
        weight_rom[9256] = 19;
        weight_rom[9257] = 9;
        weight_rom[9258] = 17;
        weight_rom[9259] = 9;
        weight_rom[9260] = 11;
        weight_rom[9261] = 17;
        weight_rom[9262] = 25;
        weight_rom[9263] = 10;
        weight_rom[9264] = 8;
        weight_rom[9265] = 9;
        weight_rom[9266] = -2;
        weight_rom[9267] = 3;
        weight_rom[9268] = -2;
        weight_rom[9269] = 0;
        weight_rom[9270] = 1;
        weight_rom[9271] = 26;
        weight_rom[9272] = 20;
        weight_rom[9273] = 21;
        weight_rom[9274] = 8;
        weight_rom[9275] = 17;
        weight_rom[9276] = 30;
        weight_rom[9277] = 34;
        weight_rom[9278] = 32;
        weight_rom[9279] = 30;
        weight_rom[9280] = 29;
        weight_rom[9281] = 25;
        weight_rom[9282] = 30;
        weight_rom[9283] = 30;
        weight_rom[9284] = 22;
        weight_rom[9285] = 8;
        weight_rom[9286] = 13;
        weight_rom[9287] = 18;
        weight_rom[9288] = 23;
        weight_rom[9289] = 5;
        weight_rom[9290] = 21;
        weight_rom[9291] = 33;
        weight_rom[9292] = 19;
        weight_rom[9293] = 8;
        weight_rom[9294] = -14;
        weight_rom[9295] = 2;
        weight_rom[9296] = -4;
        weight_rom[9297] = 4;
        weight_rom[9298] = 3;
        weight_rom[9299] = 17;
        weight_rom[9300] = 4;
        weight_rom[9301] = -10;
        weight_rom[9302] = 4;
        weight_rom[9303] = 9;
        weight_rom[9304] = 14;
        weight_rom[9305] = 26;
        weight_rom[9306] = 12;
        weight_rom[9307] = 28;
        weight_rom[9308] = 36;
        weight_rom[9309] = 34;
        weight_rom[9310] = 38;
        weight_rom[9311] = 40;
        weight_rom[9312] = 35;
        weight_rom[9313] = 31;
        weight_rom[9314] = 32;
        weight_rom[9315] = 16;
        weight_rom[9316] = 1;
        weight_rom[9317] = 9;
        weight_rom[9318] = 6;
        weight_rom[9319] = 10;
        weight_rom[9320] = 24;
        weight_rom[9321] = 19;
        weight_rom[9322] = 1;
        weight_rom[9323] = 1;
        weight_rom[9324] = -2;
        weight_rom[9325] = -2;
        weight_rom[9326] = 2;
        weight_rom[9327] = 10;
        weight_rom[9328] = 0;
        weight_rom[9329] = -8;
        weight_rom[9330] = 16;
        weight_rom[9331] = 1;
        weight_rom[9332] = 14;
        weight_rom[9333] = 9;
        weight_rom[9334] = 20;
        weight_rom[9335] = 14;
        weight_rom[9336] = 33;
        weight_rom[9337] = 26;
        weight_rom[9338] = 13;
        weight_rom[9339] = 30;
        weight_rom[9340] = 31;
        weight_rom[9341] = 40;
        weight_rom[9342] = 20;
        weight_rom[9343] = 22;
        weight_rom[9344] = -3;
        weight_rom[9345] = 7;
        weight_rom[9346] = 30;
        weight_rom[9347] = 14;
        weight_rom[9348] = 17;
        weight_rom[9349] = 4;
        weight_rom[9350] = 4;
        weight_rom[9351] = -4;
        weight_rom[9352] = -1;
        weight_rom[9353] = 0;
        weight_rom[9354] = 2;
        weight_rom[9355] = -2;
        weight_rom[9356] = -11;
        weight_rom[9357] = -23;
        weight_rom[9358] = -20;
        weight_rom[9359] = -17;
        weight_rom[9360] = -18;
        weight_rom[9361] = 1;
        weight_rom[9362] = 1;
        weight_rom[9363] = 9;
        weight_rom[9364] = 15;
        weight_rom[9365] = 12;
        weight_rom[9366] = -5;
        weight_rom[9367] = 11;
        weight_rom[9368] = 11;
        weight_rom[9369] = -2;
        weight_rom[9370] = -3;
        weight_rom[9371] = 10;
        weight_rom[9372] = 3;
        weight_rom[9373] = 7;
        weight_rom[9374] = 9;
        weight_rom[9375] = -1;
        weight_rom[9376] = -2;
        weight_rom[9377] = 1;
        weight_rom[9378] = 0;
        weight_rom[9379] = -1;
        weight_rom[9380] = -4;
        weight_rom[9381] = 4;
        weight_rom[9382] = 1;
        weight_rom[9383] = 1;
        weight_rom[9384] = 1;
        weight_rom[9385] = 2;
        weight_rom[9386] = 0;
        weight_rom[9387] = 9;
        weight_rom[9388] = 11;
        weight_rom[9389] = -8;
        weight_rom[9390] = 5;
        weight_rom[9391] = 15;
        weight_rom[9392] = 10;
        weight_rom[9393] = 3;
        weight_rom[9394] = -1;
        weight_rom[9395] = -9;
        weight_rom[9396] = -9;
        weight_rom[9397] = 0;
        weight_rom[9398] = -8;
        weight_rom[9399] = 0;
        weight_rom[9400] = 1;
        weight_rom[9401] = 0;
        weight_rom[9402] = -6;
        weight_rom[9403] = 2;
        weight_rom[9404] = -2;
        weight_rom[9405] = -1;
        weight_rom[9406] = -3;
        weight_rom[9407] = -1;
        weight_rom[9408] = -4;
        weight_rom[9409] = 2;
        weight_rom[9410] = 1;
        weight_rom[9411] = 4;
        weight_rom[9412] = -3;
        weight_rom[9413] = -1;
        weight_rom[9414] = -1;
        weight_rom[9415] = 4;
        weight_rom[9416] = -4;
        weight_rom[9417] = 0;
        weight_rom[9418] = 0;
        weight_rom[9419] = 2;
        weight_rom[9420] = 4;
        weight_rom[9421] = -3;
        weight_rom[9422] = -2;
        weight_rom[9423] = -3;
        weight_rom[9424] = 0;
        weight_rom[9425] = -4;
        weight_rom[9426] = 0;
        weight_rom[9427] = 0;
        weight_rom[9428] = 4;
        weight_rom[9429] = 0;
        weight_rom[9430] = -4;
        weight_rom[9431] = -5;
        weight_rom[9432] = 0;
        weight_rom[9433] = 0;
        weight_rom[9434] = 2;
        weight_rom[9435] = -2;
        weight_rom[9436] = -2;
        weight_rom[9437] = 3;
        weight_rom[9438] = 0;
        weight_rom[9439] = -1;
        weight_rom[9440] = 4;
        weight_rom[9441] = 0;
        weight_rom[9442] = -13;
        weight_rom[9443] = -23;
        weight_rom[9444] = -18;
        weight_rom[9445] = -8;
        weight_rom[9446] = -22;
        weight_rom[9447] = 1;
        weight_rom[9448] = -21;
        weight_rom[9449] = -25;
        weight_rom[9450] = -1;
        weight_rom[9451] = -33;
        weight_rom[9452] = -37;
        weight_rom[9453] = -20;
        weight_rom[9454] = -21;
        weight_rom[9455] = -28;
        weight_rom[9456] = -21;
        weight_rom[9457] = -18;
        weight_rom[9458] = -18;
        weight_rom[9459] = -10;
        weight_rom[9460] = 3;
        weight_rom[9461] = 3;
        weight_rom[9462] = -4;
        weight_rom[9463] = -2;
        weight_rom[9464] = -3;
        weight_rom[9465] = -2;
        weight_rom[9466] = 0;
        weight_rom[9467] = -1;
        weight_rom[9468] = -9;
        weight_rom[9469] = 2;
        weight_rom[9470] = -22;
        weight_rom[9471] = -35;
        weight_rom[9472] = -38;
        weight_rom[9473] = -40;
        weight_rom[9474] = -49;
        weight_rom[9475] = -44;
        weight_rom[9476] = -54;
        weight_rom[9477] = -30;
        weight_rom[9478] = -28;
        weight_rom[9479] = -26;
        weight_rom[9480] = -39;
        weight_rom[9481] = -42;
        weight_rom[9482] = -38;
        weight_rom[9483] = -21;
        weight_rom[9484] = -33;
        weight_rom[9485] = -36;
        weight_rom[9486] = -22;
        weight_rom[9487] = -29;
        weight_rom[9488] = -26;
        weight_rom[9489] = -9;
        weight_rom[9490] = 2;
        weight_rom[9491] = -4;
        weight_rom[9492] = -3;
        weight_rom[9493] = 4;
        weight_rom[9494] = -12;
        weight_rom[9495] = -1;
        weight_rom[9496] = 0;
        weight_rom[9497] = -17;
        weight_rom[9498] = -36;
        weight_rom[9499] = -35;
        weight_rom[9500] = -45;
        weight_rom[9501] = -70;
        weight_rom[9502] = -55;
        weight_rom[9503] = -46;
        weight_rom[9504] = -50;
        weight_rom[9505] = -60;
        weight_rom[9506] = -23;
        weight_rom[9507] = -40;
        weight_rom[9508] = -15;
        weight_rom[9509] = -10;
        weight_rom[9510] = -30;
        weight_rom[9511] = -23;
        weight_rom[9512] = -27;
        weight_rom[9513] = -20;
        weight_rom[9514] = -28;
        weight_rom[9515] = -20;
        weight_rom[9516] = -26;
        weight_rom[9517] = 18;
        weight_rom[9518] = 4;
        weight_rom[9519] = 2;
        weight_rom[9520] = 0;
        weight_rom[9521] = 2;
        weight_rom[9522] = -1;
        weight_rom[9523] = -4;
        weight_rom[9524] = -9;
        weight_rom[9525] = -26;
        weight_rom[9526] = -27;
        weight_rom[9527] = -12;
        weight_rom[9528] = -26;
        weight_rom[9529] = -24;
        weight_rom[9530] = -37;
        weight_rom[9531] = -15;
        weight_rom[9532] = -22;
        weight_rom[9533] = -22;
        weight_rom[9534] = -26;
        weight_rom[9535] = -15;
        weight_rom[9536] = -9;
        weight_rom[9537] = -6;
        weight_rom[9538] = -21;
        weight_rom[9539] = -15;
        weight_rom[9540] = -3;
        weight_rom[9541] = 19;
        weight_rom[9542] = 25;
        weight_rom[9543] = 16;
        weight_rom[9544] = 37;
        weight_rom[9545] = 6;
        weight_rom[9546] = 8;
        weight_rom[9547] = 2;
        weight_rom[9548] = 3;
        weight_rom[9549] = -2;
        weight_rom[9550] = -1;
        weight_rom[9551] = -8;
        weight_rom[9552] = -24;
        weight_rom[9553] = -13;
        weight_rom[9554] = -14;
        weight_rom[9555] = -7;
        weight_rom[9556] = -10;
        weight_rom[9557] = 2;
        weight_rom[9558] = 3;
        weight_rom[9559] = 8;
        weight_rom[9560] = 3;
        weight_rom[9561] = -10;
        weight_rom[9562] = 1;
        weight_rom[9563] = -1;
        weight_rom[9564] = 3;
        weight_rom[9565] = 8;
        weight_rom[9566] = 1;
        weight_rom[9567] = -11;
        weight_rom[9568] = 3;
        weight_rom[9569] = 2;
        weight_rom[9570] = 17;
        weight_rom[9571] = 29;
        weight_rom[9572] = 10;
        weight_rom[9573] = 0;
        weight_rom[9574] = -13;
        weight_rom[9575] = -4;
        weight_rom[9576] = 1;
        weight_rom[9577] = 1;
        weight_rom[9578] = -1;
        weight_rom[9579] = -21;
        weight_rom[9580] = -4;
        weight_rom[9581] = 0;
        weight_rom[9582] = -6;
        weight_rom[9583] = 1;
        weight_rom[9584] = -1;
        weight_rom[9585] = 2;
        weight_rom[9586] = 6;
        weight_rom[9587] = -1;
        weight_rom[9588] = 0;
        weight_rom[9589] = -9;
        weight_rom[9590] = -5;
        weight_rom[9591] = -14;
        weight_rom[9592] = -9;
        weight_rom[9593] = 8;
        weight_rom[9594] = 12;
        weight_rom[9595] = 14;
        weight_rom[9596] = 15;
        weight_rom[9597] = 25;
        weight_rom[9598] = 31;
        weight_rom[9599] = 30;
        weight_rom[9600] = 25;
        weight_rom[9601] = 11;
        weight_rom[9602] = 21;
        weight_rom[9603] = -24;
        weight_rom[9604] = 0;
        weight_rom[9605] = -17;
        weight_rom[9606] = 6;
        weight_rom[9607] = -15;
        weight_rom[9608] = -23;
        weight_rom[9609] = 7;
        weight_rom[9610] = -1;
        weight_rom[9611] = 7;
        weight_rom[9612] = 0;
        weight_rom[9613] = 6;
        weight_rom[9614] = 0;
        weight_rom[9615] = 3;
        weight_rom[9616] = -10;
        weight_rom[9617] = 0;
        weight_rom[9618] = -16;
        weight_rom[9619] = -10;
        weight_rom[9620] = 3;
        weight_rom[9621] = 16;
        weight_rom[9622] = 16;
        weight_rom[9623] = 23;
        weight_rom[9624] = 28;
        weight_rom[9625] = 26;
        weight_rom[9626] = 33;
        weight_rom[9627] = 43;
        weight_rom[9628] = 17;
        weight_rom[9629] = 26;
        weight_rom[9630] = 14;
        weight_rom[9631] = 3;
        weight_rom[9632] = -1;
        weight_rom[9633] = -14;
        weight_rom[9634] = 7;
        weight_rom[9635] = -23;
        weight_rom[9636] = -26;
        weight_rom[9637] = 5;
        weight_rom[9638] = -4;
        weight_rom[9639] = -19;
        weight_rom[9640] = 5;
        weight_rom[9641] = 5;
        weight_rom[9642] = 0;
        weight_rom[9643] = 1;
        weight_rom[9644] = -14;
        weight_rom[9645] = -13;
        weight_rom[9646] = -18;
        weight_rom[9647] = -1;
        weight_rom[9648] = 10;
        weight_rom[9649] = 18;
        weight_rom[9650] = 30;
        weight_rom[9651] = 24;
        weight_rom[9652] = 24;
        weight_rom[9653] = 22;
        weight_rom[9654] = 20;
        weight_rom[9655] = 34;
        weight_rom[9656] = 47;
        weight_rom[9657] = 37;
        weight_rom[9658] = -1;
        weight_rom[9659] = -14;
        weight_rom[9660] = -6;
        weight_rom[9661] = -13;
        weight_rom[9662] = -2;
        weight_rom[9663] = -19;
        weight_rom[9664] = -26;
        weight_rom[9665] = -5;
        weight_rom[9666] = -7;
        weight_rom[9667] = -13;
        weight_rom[9668] = -1;
        weight_rom[9669] = 1;
        weight_rom[9670] = 11;
        weight_rom[9671] = 0;
        weight_rom[9672] = 4;
        weight_rom[9673] = 1;
        weight_rom[9674] = -22;
        weight_rom[9675] = -10;
        weight_rom[9676] = 16;
        weight_rom[9677] = 23;
        weight_rom[9678] = 34;
        weight_rom[9679] = 23;
        weight_rom[9680] = 20;
        weight_rom[9681] = 22;
        weight_rom[9682] = 13;
        weight_rom[9683] = 27;
        weight_rom[9684] = 37;
        weight_rom[9685] = 24;
        weight_rom[9686] = 2;
        weight_rom[9687] = -3;
        weight_rom[9688] = -12;
        weight_rom[9689] = -6;
        weight_rom[9690] = -4;
        weight_rom[9691] = -35;
        weight_rom[9692] = -21;
        weight_rom[9693] = -8;
        weight_rom[9694] = -13;
        weight_rom[9695] = -5;
        weight_rom[9696] = 12;
        weight_rom[9697] = 14;
        weight_rom[9698] = 14;
        weight_rom[9699] = 15;
        weight_rom[9700] = 9;
        weight_rom[9701] = -16;
        weight_rom[9702] = -31;
        weight_rom[9703] = -15;
        weight_rom[9704] = 5;
        weight_rom[9705] = 22;
        weight_rom[9706] = 13;
        weight_rom[9707] = 14;
        weight_rom[9708] = 7;
        weight_rom[9709] = 7;
        weight_rom[9710] = 4;
        weight_rom[9711] = -7;
        weight_rom[9712] = 21;
        weight_rom[9713] = 36;
        weight_rom[9714] = -12;
        weight_rom[9715] = 6;
        weight_rom[9716] = 6;
        weight_rom[9717] = -16;
        weight_rom[9718] = -32;
        weight_rom[9719] = -23;
        weight_rom[9720] = -38;
        weight_rom[9721] = -14;
        weight_rom[9722] = 13;
        weight_rom[9723] = 5;
        weight_rom[9724] = 18;
        weight_rom[9725] = 18;
        weight_rom[9726] = 19;
        weight_rom[9727] = 10;
        weight_rom[9728] = 10;
        weight_rom[9729] = -24;
        weight_rom[9730] = -52;
        weight_rom[9731] = -20;
        weight_rom[9732] = 0;
        weight_rom[9733] = 9;
        weight_rom[9734] = 6;
        weight_rom[9735] = -4;
        weight_rom[9736] = -8;
        weight_rom[9737] = -4;
        weight_rom[9738] = -15;
        weight_rom[9739] = -23;
        weight_rom[9740] = -18;
        weight_rom[9741] = 4;
        weight_rom[9742] = 20;
        weight_rom[9743] = -13;
        weight_rom[9744] = 6;
        weight_rom[9745] = -8;
        weight_rom[9746] = -21;
        weight_rom[9747] = -29;
        weight_rom[9748] = -23;
        weight_rom[9749] = -10;
        weight_rom[9750] = 24;
        weight_rom[9751] = 17;
        weight_rom[9752] = 25;
        weight_rom[9753] = 19;
        weight_rom[9754] = 27;
        weight_rom[9755] = 27;
        weight_rom[9756] = 15;
        weight_rom[9757] = -10;
        weight_rom[9758] = -40;
        weight_rom[9759] = -25;
        weight_rom[9760] = -8;
        weight_rom[9761] = -3;
        weight_rom[9762] = -5;
        weight_rom[9763] = 1;
        weight_rom[9764] = -7;
        weight_rom[9765] = -5;
        weight_rom[9766] = -13;
        weight_rom[9767] = -24;
        weight_rom[9768] = -27;
        weight_rom[9769] = -19;
        weight_rom[9770] = -12;
        weight_rom[9771] = -12;
        weight_rom[9772] = -4;
        weight_rom[9773] = 2;
        weight_rom[9774] = -26;
        weight_rom[9775] = -34;
        weight_rom[9776] = 4;
        weight_rom[9777] = 16;
        weight_rom[9778] = 30;
        weight_rom[9779] = 44;
        weight_rom[9780] = 31;
        weight_rom[9781] = 26;
        weight_rom[9782] = 30;
        weight_rom[9783] = 27;
        weight_rom[9784] = 11;
        weight_rom[9785] = -14;
        weight_rom[9786] = -26;
        weight_rom[9787] = -23;
        weight_rom[9788] = -8;
        weight_rom[9789] = 6;
        weight_rom[9790] = 6;
        weight_rom[9791] = 0;
        weight_rom[9792] = 12;
        weight_rom[9793] = 3;
        weight_rom[9794] = -2;
        weight_rom[9795] = -14;
        weight_rom[9796] = -25;
        weight_rom[9797] = -4;
        weight_rom[9798] = -16;
        weight_rom[9799] = -16;
        weight_rom[9800] = -3;
        weight_rom[9801] = -7;
        weight_rom[9802] = -3;
        weight_rom[9803] = -17;
        weight_rom[9804] = 35;
        weight_rom[9805] = 24;
        weight_rom[9806] = 29;
        weight_rom[9807] = 41;
        weight_rom[9808] = 25;
        weight_rom[9809] = 30;
        weight_rom[9810] = 22;
        weight_rom[9811] = 21;
        weight_rom[9812] = 11;
        weight_rom[9813] = -5;
        weight_rom[9814] = -15;
        weight_rom[9815] = -19;
        weight_rom[9816] = -2;
        weight_rom[9817] = 19;
        weight_rom[9818] = 9;
        weight_rom[9819] = 4;
        weight_rom[9820] = -2;
        weight_rom[9821] = -4;
        weight_rom[9822] = 3;
        weight_rom[9823] = -3;
        weight_rom[9824] = 12;
        weight_rom[9825] = -23;
        weight_rom[9826] = -33;
        weight_rom[9827] = 4;
        weight_rom[9828] = 4;
        weight_rom[9829] = -8;
        weight_rom[9830] = -7;
        weight_rom[9831] = 4;
        weight_rom[9832] = 27;
        weight_rom[9833] = 24;
        weight_rom[9834] = 18;
        weight_rom[9835] = 29;
        weight_rom[9836] = 38;
        weight_rom[9837] = 27;
        weight_rom[9838] = 25;
        weight_rom[9839] = 22;
        weight_rom[9840] = 10;
        weight_rom[9841] = -20;
        weight_rom[9842] = -21;
        weight_rom[9843] = -7;
        weight_rom[9844] = 12;
        weight_rom[9845] = 20;
        weight_rom[9846] = 16;
        weight_rom[9847] = 4;
        weight_rom[9848] = -3;
        weight_rom[9849] = -12;
        weight_rom[9850] = -6;
        weight_rom[9851] = 2;
        weight_rom[9852] = -17;
        weight_rom[9853] = -29;
        weight_rom[9854] = -1;
        weight_rom[9855] = -18;
        weight_rom[9856] = -1;
        weight_rom[9857] = -1;
        weight_rom[9858] = -23;
        weight_rom[9859] = -19;
        weight_rom[9860] = -17;
        weight_rom[9861] = 11;
        weight_rom[9862] = 16;
        weight_rom[9863] = 13;
        weight_rom[9864] = 27;
        weight_rom[9865] = 6;
        weight_rom[9866] = 9;
        weight_rom[9867] = 7;
        weight_rom[9868] = 2;
        weight_rom[9869] = -7;
        weight_rom[9870] = -5;
        weight_rom[9871] = 6;
        weight_rom[9872] = 18;
        weight_rom[9873] = 16;
        weight_rom[9874] = 13;
        weight_rom[9875] = 0;
        weight_rom[9876] = 2;
        weight_rom[9877] = -3;
        weight_rom[9878] = -5;
        weight_rom[9879] = -3;
        weight_rom[9880] = -8;
        weight_rom[9881] = -34;
        weight_rom[9882] = -20;
        weight_rom[9883] = -18;
        weight_rom[9884] = -3;
        weight_rom[9885] = -1;
        weight_rom[9886] = 0;
        weight_rom[9887] = -28;
        weight_rom[9888] = -12;
        weight_rom[9889] = 8;
        weight_rom[9890] = 11;
        weight_rom[9891] = 2;
        weight_rom[9892] = 12;
        weight_rom[9893] = 1;
        weight_rom[9894] = -2;
        weight_rom[9895] = -12;
        weight_rom[9896] = -6;
        weight_rom[9897] = -6;
        weight_rom[9898] = 3;
        weight_rom[9899] = 22;
        weight_rom[9900] = 20;
        weight_rom[9901] = 20;
        weight_rom[9902] = 9;
        weight_rom[9903] = -2;
        weight_rom[9904] = -1;
        weight_rom[9905] = -2;
        weight_rom[9906] = -11;
        weight_rom[9907] = -13;
        weight_rom[9908] = -9;
        weight_rom[9909] = -23;
        weight_rom[9910] = -21;
        weight_rom[9911] = -2;
        weight_rom[9912] = 4;
        weight_rom[9913] = -2;
        weight_rom[9914] = -11;
        weight_rom[9915] = -17;
        weight_rom[9916] = 7;
        weight_rom[9917] = 12;
        weight_rom[9918] = 15;
        weight_rom[9919] = 2;
        weight_rom[9920] = 6;
        weight_rom[9921] = -12;
        weight_rom[9922] = -9;
        weight_rom[9923] = -1;
        weight_rom[9924] = -5;
        weight_rom[9925] = -5;
        weight_rom[9926] = 6;
        weight_rom[9927] = 9;
        weight_rom[9928] = 9;
        weight_rom[9929] = -2;
        weight_rom[9930] = -12;
        weight_rom[9931] = -4;
        weight_rom[9932] = 6;
        weight_rom[9933] = -1;
        weight_rom[9934] = -17;
        weight_rom[9935] = -24;
        weight_rom[9936] = -23;
        weight_rom[9937] = -35;
        weight_rom[9938] = -17;
        weight_rom[9939] = -6;
        weight_rom[9940] = 2;
        weight_rom[9941] = -8;
        weight_rom[9942] = 3;
        weight_rom[9943] = -5;
        weight_rom[9944] = 12;
        weight_rom[9945] = 18;
        weight_rom[9946] = 9;
        weight_rom[9947] = 0;
        weight_rom[9948] = -11;
        weight_rom[9949] = -14;
        weight_rom[9950] = -10;
        weight_rom[9951] = 1;
        weight_rom[9952] = -10;
        weight_rom[9953] = -2;
        weight_rom[9954] = -11;
        weight_rom[9955] = -4;
        weight_rom[9956] = -6;
        weight_rom[9957] = -10;
        weight_rom[9958] = -5;
        weight_rom[9959] = -7;
        weight_rom[9960] = -4;
        weight_rom[9961] = -11;
        weight_rom[9962] = -28;
        weight_rom[9963] = -23;
        weight_rom[9964] = 1;
        weight_rom[9965] = 3;
        weight_rom[9966] = -1;
        weight_rom[9967] = 4;
        weight_rom[9968] = -3;
        weight_rom[9969] = 5;
        weight_rom[9970] = -3;
        weight_rom[9971] = -16;
        weight_rom[9972] = -7;
        weight_rom[9973] = -2;
        weight_rom[9974] = 1;
        weight_rom[9975] = -22;
        weight_rom[9976] = -11;
        weight_rom[9977] = -10;
        weight_rom[9978] = -10;
        weight_rom[9979] = 5;
        weight_rom[9980] = -7;
        weight_rom[9981] = -8;
        weight_rom[9982] = -11;
        weight_rom[9983] = -6;
        weight_rom[9984] = 1;
        weight_rom[9985] = 2;
        weight_rom[9986] = 2;
        weight_rom[9987] = -14;
        weight_rom[9988] = -12;
        weight_rom[9989] = -12;
        weight_rom[9990] = 4;
        weight_rom[9991] = -15;
        weight_rom[9992] = -6;
        weight_rom[9993] = -6;
        weight_rom[9994] = -13;
        weight_rom[9995] = 1;
        weight_rom[9996] = 4;
        weight_rom[9997] = -8;
        weight_rom[9998] = -27;
        weight_rom[9999] = -16;
        weight_rom[10000] = -5;
        weight_rom[10001] = -1;
        weight_rom[10002] = -13;
        weight_rom[10003] = -20;
        weight_rom[10004] = -17;
        weight_rom[10005] = 2;
        weight_rom[10006] = -15;
        weight_rom[10007] = -11;
        weight_rom[10008] = -12;
        weight_rom[10009] = -20;
        weight_rom[10010] = -16;
        weight_rom[10011] = -5;
        weight_rom[10012] = -8;
        weight_rom[10013] = -4;
        weight_rom[10014] = -3;
        weight_rom[10015] = -3;
        weight_rom[10016] = 5;
        weight_rom[10017] = 10;
        weight_rom[10018] = 4;
        weight_rom[10019] = 10;
        weight_rom[10020] = -4;
        weight_rom[10021] = -11;
        weight_rom[10022] = -10;
        weight_rom[10023] = 2;
        weight_rom[10024] = 0;
        weight_rom[10025] = 1;
        weight_rom[10026] = -25;
        weight_rom[10027] = -29;
        weight_rom[10028] = -11;
        weight_rom[10029] = -20;
        weight_rom[10030] = -1;
        weight_rom[10031] = -8;
        weight_rom[10032] = 8;
        weight_rom[10033] = -2;
        weight_rom[10034] = 2;
        weight_rom[10035] = 3;
        weight_rom[10036] = -2;
        weight_rom[10037] = 0;
        weight_rom[10038] = -5;
        weight_rom[10039] = -11;
        weight_rom[10040] = 3;
        weight_rom[10041] = 3;
        weight_rom[10042] = -4;
        weight_rom[10043] = 6;
        weight_rom[10044] = 9;
        weight_rom[10045] = 26;
        weight_rom[10046] = 18;
        weight_rom[10047] = 15;
        weight_rom[10048] = 3;
        weight_rom[10049] = 4;
        weight_rom[10050] = -1;
        weight_rom[10051] = -2;
        weight_rom[10052] = -4;
        weight_rom[10053] = 4;
        weight_rom[10054] = -21;
        weight_rom[10055] = -10;
        weight_rom[10056] = -34;
        weight_rom[10057] = -4;
        weight_rom[10058] = -1;
        weight_rom[10059] = 2;
        weight_rom[10060] = 11;
        weight_rom[10061] = 11;
        weight_rom[10062] = 18;
        weight_rom[10063] = 18;
        weight_rom[10064] = 13;
        weight_rom[10065] = 10;
        weight_rom[10066] = 16;
        weight_rom[10067] = 3;
        weight_rom[10068] = 24;
        weight_rom[10069] = 22;
        weight_rom[10070] = 16;
        weight_rom[10071] = 6;
        weight_rom[10072] = 17;
        weight_rom[10073] = 21;
        weight_rom[10074] = 3;
        weight_rom[10075] = -6;
        weight_rom[10076] = -2;
        weight_rom[10077] = 17;
        weight_rom[10078] = 3;
        weight_rom[10079] = 3;
        weight_rom[10080] = 0;
        weight_rom[10081] = -1;
        weight_rom[10082] = -6;
        weight_rom[10083] = -8;
        weight_rom[10084] = -14;
        weight_rom[10085] = 7;
        weight_rom[10086] = 16;
        weight_rom[10087] = 6;
        weight_rom[10088] = 8;
        weight_rom[10089] = 10;
        weight_rom[10090] = 11;
        weight_rom[10091] = 8;
        weight_rom[10092] = 10;
        weight_rom[10093] = 3;
        weight_rom[10094] = 1;
        weight_rom[10095] = 10;
        weight_rom[10096] = -2;
        weight_rom[10097] = 12;
        weight_rom[10098] = 5;
        weight_rom[10099] = 2;
        weight_rom[10100] = 10;
        weight_rom[10101] = -5;
        weight_rom[10102] = 31;
        weight_rom[10103] = 13;
        weight_rom[10104] = -1;
        weight_rom[10105] = -24;
        weight_rom[10106] = 1;
        weight_rom[10107] = 4;
        weight_rom[10108] = 3;
        weight_rom[10109] = 1;
        weight_rom[10110] = 2;
        weight_rom[10111] = 10;
        weight_rom[10112] = 15;
        weight_rom[10113] = 10;
        weight_rom[10114] = -5;
        weight_rom[10115] = -20;
        weight_rom[10116] = -32;
        weight_rom[10117] = -23;
        weight_rom[10118] = -20;
        weight_rom[10119] = -24;
        weight_rom[10120] = -31;
        weight_rom[10121] = -13;
        weight_rom[10122] = -17;
        weight_rom[10123] = -17;
        weight_rom[10124] = -18;
        weight_rom[10125] = -26;
        weight_rom[10126] = -18;
        weight_rom[10127] = -20;
        weight_rom[10128] = -16;
        weight_rom[10129] = -10;
        weight_rom[10130] = 5;
        weight_rom[10131] = 5;
        weight_rom[10132] = -6;
        weight_rom[10133] = 4;
        weight_rom[10134] = -4;
        weight_rom[10135] = -4;
        weight_rom[10136] = -1;
        weight_rom[10137] = 2;
        weight_rom[10138] = 0;
        weight_rom[10139] = 0;
        weight_rom[10140] = 13;
        weight_rom[10141] = 16;
        weight_rom[10142] = -1;
        weight_rom[10143] = -28;
        weight_rom[10144] = -28;
        weight_rom[10145] = -42;
        weight_rom[10146] = -23;
        weight_rom[10147] = -26;
        weight_rom[10148] = -10;
        weight_rom[10149] = -37;
        weight_rom[10150] = -35;
        weight_rom[10151] = -20;
        weight_rom[10152] = -31;
        weight_rom[10153] = -39;
        weight_rom[10154] = -30;
        weight_rom[10155] = -38;
        weight_rom[10156] = -11;
        weight_rom[10157] = -14;
        weight_rom[10158] = -29;
        weight_rom[10159] = -10;
        weight_rom[10160] = -3;
        weight_rom[10161] = -4;
        weight_rom[10162] = 4;
        weight_rom[10163] = 4;
        weight_rom[10164] = 2;
        weight_rom[10165] = -2;
        weight_rom[10166] = -2;
        weight_rom[10167] = 4;
        weight_rom[10168] = -4;
        weight_rom[10169] = -23;
        weight_rom[10170] = -11;
        weight_rom[10171] = -23;
        weight_rom[10172] = -27;
        weight_rom[10173] = -13;
        weight_rom[10174] = -24;
        weight_rom[10175] = -10;
        weight_rom[10176] = -18;
        weight_rom[10177] = -21;
        weight_rom[10178] = -31;
        weight_rom[10179] = -16;
        weight_rom[10180] = -10;
        weight_rom[10181] = -24;
        weight_rom[10182] = -21;
        weight_rom[10183] = -15;
        weight_rom[10184] = -9;
        weight_rom[10185] = -10;
        weight_rom[10186] = -19;
        weight_rom[10187] = -4;
        weight_rom[10188] = -1;
        weight_rom[10189] = 0;
        weight_rom[10190] = 1;
        weight_rom[10191] = -1;
        weight_rom[10192] = 1;
        weight_rom[10193] = 0;
        weight_rom[10194] = 4;
        weight_rom[10195] = -2;
        weight_rom[10196] = -3;
        weight_rom[10197] = -4;
        weight_rom[10198] = 0;
        weight_rom[10199] = 2;
        weight_rom[10200] = 1;
        weight_rom[10201] = -1;
        weight_rom[10202] = -3;
        weight_rom[10203] = -1;
        weight_rom[10204] = 4;
        weight_rom[10205] = 7;
        weight_rom[10206] = 6;
        weight_rom[10207] = 1;
        weight_rom[10208] = 0;
        weight_rom[10209] = -1;
        weight_rom[10210] = 4;
        weight_rom[10211] = 4;
        weight_rom[10212] = -4;
        weight_rom[10213] = 2;
        weight_rom[10214] = -3;
        weight_rom[10215] = 1;
        weight_rom[10216] = 4;
        weight_rom[10217] = -1;
        weight_rom[10218] = 0;
        weight_rom[10219] = 1;
        weight_rom[10220] = -3;
        weight_rom[10221] = 3;
        weight_rom[10222] = -3;
        weight_rom[10223] = 2;
        weight_rom[10224] = 2;
        weight_rom[10225] = -2;
        weight_rom[10226] = 20;
        weight_rom[10227] = 25;
        weight_rom[10228] = 17;
        weight_rom[10229] = 12;
        weight_rom[10230] = 12;
        weight_rom[10231] = 15;
        weight_rom[10232] = 19;
        weight_rom[10233] = 22;
        weight_rom[10234] = -2;
        weight_rom[10235] = 3;
        weight_rom[10236] = 35;
        weight_rom[10237] = 12;
        weight_rom[10238] = 10;
        weight_rom[10239] = 16;
        weight_rom[10240] = 13;
        weight_rom[10241] = 11;
        weight_rom[10242] = 16;
        weight_rom[10243] = 10;
        weight_rom[10244] = 0;
        weight_rom[10245] = -5;
        weight_rom[10246] = -2;
        weight_rom[10247] = -3;
        weight_rom[10248] = 3;
        weight_rom[10249] = 3;
        weight_rom[10250] = -1;
        weight_rom[10251] = 3;
        weight_rom[10252] = 2;
        weight_rom[10253] = -1;
        weight_rom[10254] = 16;
        weight_rom[10255] = 26;
        weight_rom[10256] = 25;
        weight_rom[10257] = 29;
        weight_rom[10258] = 30;
        weight_rom[10259] = 27;
        weight_rom[10260] = 25;
        weight_rom[10261] = -9;
        weight_rom[10262] = 1;
        weight_rom[10263] = -17;
        weight_rom[10264] = 10;
        weight_rom[10265] = 11;
        weight_rom[10266] = 40;
        weight_rom[10267] = 9;
        weight_rom[10268] = 26;
        weight_rom[10269] = 16;
        weight_rom[10270] = 15;
        weight_rom[10271] = 9;
        weight_rom[10272] = -1;
        weight_rom[10273] = -11;
        weight_rom[10274] = 0;
        weight_rom[10275] = -3;
        weight_rom[10276] = 1;
        weight_rom[10277] = 2;
        weight_rom[10278] = 8;
        weight_rom[10279] = 0;
        weight_rom[10280] = 2;
        weight_rom[10281] = 18;
        weight_rom[10282] = 29;
        weight_rom[10283] = 34;
        weight_rom[10284] = 40;
        weight_rom[10285] = 23;
        weight_rom[10286] = 34;
        weight_rom[10287] = 57;
        weight_rom[10288] = 39;
        weight_rom[10289] = 17;
        weight_rom[10290] = 24;
        weight_rom[10291] = 16;
        weight_rom[10292] = 13;
        weight_rom[10293] = 37;
        weight_rom[10294] = 41;
        weight_rom[10295] = 45;
        weight_rom[10296] = 48;
        weight_rom[10297] = 33;
        weight_rom[10298] = 39;
        weight_rom[10299] = 31;
        weight_rom[10300] = 28;
        weight_rom[10301] = 3;
        weight_rom[10302] = 3;
        weight_rom[10303] = 1;
        weight_rom[10304] = 0;
        weight_rom[10305] = -3;
        weight_rom[10306] = -14;
        weight_rom[10307] = 0;
        weight_rom[10308] = 9;
        weight_rom[10309] = 11;
        weight_rom[10310] = 8;
        weight_rom[10311] = 30;
        weight_rom[10312] = 18;
        weight_rom[10313] = 39;
        weight_rom[10314] = 49;
        weight_rom[10315] = 39;
        weight_rom[10316] = 38;
        weight_rom[10317] = 19;
        weight_rom[10318] = 35;
        weight_rom[10319] = 31;
        weight_rom[10320] = 39;
        weight_rom[10321] = 39;
        weight_rom[10322] = 33;
        weight_rom[10323] = 25;
        weight_rom[10324] = 15;
        weight_rom[10325] = 24;
        weight_rom[10326] = 21;
        weight_rom[10327] = 16;
        weight_rom[10328] = 44;
        weight_rom[10329] = 24;
        weight_rom[10330] = 14;
        weight_rom[10331] = -1;
        weight_rom[10332] = 4;
        weight_rom[10333] = 3;
        weight_rom[10334] = 3;
        weight_rom[10335] = 0;
        weight_rom[10336] = 8;
        weight_rom[10337] = -19;
        weight_rom[10338] = -9;
        weight_rom[10339] = 7;
        weight_rom[10340] = -5;
        weight_rom[10341] = 6;
        weight_rom[10342] = 13;
        weight_rom[10343] = 13;
        weight_rom[10344] = 9;
        weight_rom[10345] = 10;
        weight_rom[10346] = 16;
        weight_rom[10347] = 29;
        weight_rom[10348] = 37;
        weight_rom[10349] = 42;
        weight_rom[10350] = 24;
        weight_rom[10351] = 25;
        weight_rom[10352] = 32;
        weight_rom[10353] = 19;
        weight_rom[10354] = 18;
        weight_rom[10355] = 22;
        weight_rom[10356] = 29;
        weight_rom[10357] = 48;
        weight_rom[10358] = 29;
        weight_rom[10359] = -2;
        weight_rom[10360] = 1;
        weight_rom[10361] = 4;
        weight_rom[10362] = 12;
        weight_rom[10363] = -1;
        weight_rom[10364] = -1;
        weight_rom[10365] = 7;
        weight_rom[10366] = 0;
        weight_rom[10367] = 6;
        weight_rom[10368] = 1;
        weight_rom[10369] = 0;
        weight_rom[10370] = -13;
        weight_rom[10371] = -19;
        weight_rom[10372] = -11;
        weight_rom[10373] = -8;
        weight_rom[10374] = -3;
        weight_rom[10375] = 4;
        weight_rom[10376] = 2;
        weight_rom[10377] = 2;
        weight_rom[10378] = -10;
        weight_rom[10379] = 6;
        weight_rom[10380] = 1;
        weight_rom[10381] = -4;
        weight_rom[10382] = 9;
        weight_rom[10383] = 36;
        weight_rom[10384] = 52;
        weight_rom[10385] = 55;
        weight_rom[10386] = 28;
        weight_rom[10387] = 14;
        weight_rom[10388] = 0;
        weight_rom[10389] = 15;
        weight_rom[10390] = -24;
        weight_rom[10391] = -12;
        weight_rom[10392] = 21;
        weight_rom[10393] = 24;
        weight_rom[10394] = 0;
        weight_rom[10395] = -6;
        weight_rom[10396] = 8;
        weight_rom[10397] = -11;
        weight_rom[10398] = -13;
        weight_rom[10399] = -14;
        weight_rom[10400] = -21;
        weight_rom[10401] = -17;
        weight_rom[10402] = -13;
        weight_rom[10403] = -14;
        weight_rom[10404] = -14;
        weight_rom[10405] = -15;
        weight_rom[10406] = -12;
        weight_rom[10407] = -11;
        weight_rom[10408] = -15;
        weight_rom[10409] = 1;
        weight_rom[10410] = 14;
        weight_rom[10411] = 19;
        weight_rom[10412] = 54;
        weight_rom[10413] = 65;
        weight_rom[10414] = 24;
        weight_rom[10415] = 4;
        weight_rom[10416] = -10;
        weight_rom[10417] = 0;
        weight_rom[10418] = 3;
        weight_rom[10419] = -4;
        weight_rom[10420] = 8;
        weight_rom[10421] = 2;
        weight_rom[10422] = 0;
        weight_rom[10423] = -1;
        weight_rom[10424] = -18;
        weight_rom[10425] = -5;
        weight_rom[10426] = -11;
        weight_rom[10427] = -13;
        weight_rom[10428] = -7;
        weight_rom[10429] = 3;
        weight_rom[10430] = -15;
        weight_rom[10431] = -12;
        weight_rom[10432] = -3;
        weight_rom[10433] = -5;
        weight_rom[10434] = -4;
        weight_rom[10435] = 7;
        weight_rom[10436] = 9;
        weight_rom[10437] = 8;
        weight_rom[10438] = 14;
        weight_rom[10439] = 24;
        weight_rom[10440] = 39;
        weight_rom[10441] = 43;
        weight_rom[10442] = 38;
        weight_rom[10443] = 9;
        weight_rom[10444] = -9;
        weight_rom[10445] = -4;
        weight_rom[10446] = -4;
        weight_rom[10447] = -13;
        weight_rom[10448] = -3;
        weight_rom[10449] = 2;
        weight_rom[10450] = -20;
        weight_rom[10451] = -15;
        weight_rom[10452] = -3;
        weight_rom[10453] = -1;
        weight_rom[10454] = -13;
        weight_rom[10455] = -5;
        weight_rom[10456] = -1;
        weight_rom[10457] = 1;
        weight_rom[10458] = -10;
        weight_rom[10459] = -13;
        weight_rom[10460] = -11;
        weight_rom[10461] = -9;
        weight_rom[10462] = 4;
        weight_rom[10463] = 14;
        weight_rom[10464] = 20;
        weight_rom[10465] = 22;
        weight_rom[10466] = 24;
        weight_rom[10467] = 36;
        weight_rom[10468] = 37;
        weight_rom[10469] = 53;
        weight_rom[10470] = 12;
        weight_rom[10471] = -16;
        weight_rom[10472] = -13;
        weight_rom[10473] = -17;
        weight_rom[10474] = -8;
        weight_rom[10475] = -2;
        weight_rom[10476] = 5;
        weight_rom[10477] = -7;
        weight_rom[10478] = -9;
        weight_rom[10479] = -4;
        weight_rom[10480] = -14;
        weight_rom[10481] = -6;
        weight_rom[10482] = -10;
        weight_rom[10483] = 3;
        weight_rom[10484] = 7;
        weight_rom[10485] = 10;
        weight_rom[10486] = -9;
        weight_rom[10487] = -11;
        weight_rom[10488] = -12;
        weight_rom[10489] = -7;
        weight_rom[10490] = 2;
        weight_rom[10491] = 2;
        weight_rom[10492] = 7;
        weight_rom[10493] = 15;
        weight_rom[10494] = 10;
        weight_rom[10495] = 14;
        weight_rom[10496] = 55;
        weight_rom[10497] = 33;
        weight_rom[10498] = 22;
        weight_rom[10499] = 15;
        weight_rom[10500] = -15;
        weight_rom[10501] = -16;
        weight_rom[10502] = -30;
        weight_rom[10503] = -15;
        weight_rom[10504] = 1;
        weight_rom[10505] = -6;
        weight_rom[10506] = -7;
        weight_rom[10507] = -18;
        weight_rom[10508] = -10;
        weight_rom[10509] = -10;
        weight_rom[10510] = -9;
        weight_rom[10511] = 6;
        weight_rom[10512] = 22;
        weight_rom[10513] = 22;
        weight_rom[10514] = 0;
        weight_rom[10515] = -18;
        weight_rom[10516] = -11;
        weight_rom[10517] = -16;
        weight_rom[10518] = -13;
        weight_rom[10519] = 2;
        weight_rom[10520] = -14;
        weight_rom[10521] = -13;
        weight_rom[10522] = -11;
        weight_rom[10523] = 12;
        weight_rom[10524] = 47;
        weight_rom[10525] = 37;
        weight_rom[10526] = 34;
        weight_rom[10527] = 8;
        weight_rom[10528] = -13;
        weight_rom[10529] = -7;
        weight_rom[10530] = -25;
        weight_rom[10531] = -18;
        weight_rom[10532] = -18;
        weight_rom[10533] = -16;
        weight_rom[10534] = -11;
        weight_rom[10535] = -6;
        weight_rom[10536] = -12;
        weight_rom[10537] = 0;
        weight_rom[10538] = 21;
        weight_rom[10539] = 26;
        weight_rom[10540] = 50;
        weight_rom[10541] = 47;
        weight_rom[10542] = 0;
        weight_rom[10543] = -11;
        weight_rom[10544] = -13;
        weight_rom[10545] = -5;
        weight_rom[10546] = -14;
        weight_rom[10547] = 7;
        weight_rom[10548] = -6;
        weight_rom[10549] = -8;
        weight_rom[10550] = -16;
        weight_rom[10551] = -6;
        weight_rom[10552] = 29;
        weight_rom[10553] = 35;
        weight_rom[10554] = 11;
        weight_rom[10555] = 4;
        weight_rom[10556] = 4;
        weight_rom[10557] = 1;
        weight_rom[10558] = -30;
        weight_rom[10559] = -23;
        weight_rom[10560] = -38;
        weight_rom[10561] = -17;
        weight_rom[10562] = -14;
        weight_rom[10563] = -16;
        weight_rom[10564] = -1;
        weight_rom[10565] = 10;
        weight_rom[10566] = 25;
        weight_rom[10567] = 47;
        weight_rom[10568] = 54;
        weight_rom[10569] = 41;
        weight_rom[10570] = 7;
        weight_rom[10571] = -4;
        weight_rom[10572] = -12;
        weight_rom[10573] = -4;
        weight_rom[10574] = 5;
        weight_rom[10575] = 6;
        weight_rom[10576] = -7;
        weight_rom[10577] = -16;
        weight_rom[10578] = -8;
        weight_rom[10579] = 16;
        weight_rom[10580] = 9;
        weight_rom[10581] = 28;
        weight_rom[10582] = 44;
        weight_rom[10583] = 25;
        weight_rom[10584] = -2;
        weight_rom[10585] = -7;
        weight_rom[10586] = -9;
        weight_rom[10587] = -22;
        weight_rom[10588] = -16;
        weight_rom[10589] = -3;
        weight_rom[10590] = -2;
        weight_rom[10591] = 0;
        weight_rom[10592] = 5;
        weight_rom[10593] = 17;
        weight_rom[10594] = 25;
        weight_rom[10595] = 40;
        weight_rom[10596] = 41;
        weight_rom[10597] = 26;
        weight_rom[10598] = 13;
        weight_rom[10599] = 6;
        weight_rom[10600] = -3;
        weight_rom[10601] = 3;
        weight_rom[10602] = 0;
        weight_rom[10603] = -4;
        weight_rom[10604] = -10;
        weight_rom[10605] = -8;
        weight_rom[10606] = -9;
        weight_rom[10607] = -13;
        weight_rom[10608] = 21;
        weight_rom[10609] = 12;
        weight_rom[10610] = 12;
        weight_rom[10611] = -3;
        weight_rom[10612] = 2;
        weight_rom[10613] = 3;
        weight_rom[10614] = 1;
        weight_rom[10615] = 0;
        weight_rom[10616] = 4;
        weight_rom[10617] = -1;
        weight_rom[10618] = -9;
        weight_rom[10619] = 5;
        weight_rom[10620] = 8;
        weight_rom[10621] = 16;
        weight_rom[10622] = 23;
        weight_rom[10623] = 22;
        weight_rom[10624] = 34;
        weight_rom[10625] = 17;
        weight_rom[10626] = 11;
        weight_rom[10627] = 9;
        weight_rom[10628] = 8;
        weight_rom[10629] = 9;
        weight_rom[10630] = 3;
        weight_rom[10631] = 10;
        weight_rom[10632] = -11;
        weight_rom[10633] = -17;
        weight_rom[10634] = -3;
        weight_rom[10635] = 8;
        weight_rom[10636] = 18;
        weight_rom[10637] = 46;
        weight_rom[10638] = 17;
        weight_rom[10639] = 7;
        weight_rom[10640] = 0;
        weight_rom[10641] = -4;
        weight_rom[10642] = 20;
        weight_rom[10643] = 22;
        weight_rom[10644] = 2;
        weight_rom[10645] = 2;
        weight_rom[10646] = 5;
        weight_rom[10647] = 10;
        weight_rom[10648] = -2;
        weight_rom[10649] = 9;
        weight_rom[10650] = 13;
        weight_rom[10651] = 20;
        weight_rom[10652] = 17;
        weight_rom[10653] = 0;
        weight_rom[10654] = 6;
        weight_rom[10655] = 6;
        weight_rom[10656] = 8;
        weight_rom[10657] = 16;
        weight_rom[10658] = 10;
        weight_rom[10659] = 7;
        weight_rom[10660] = -2;
        weight_rom[10661] = 15;
        weight_rom[10662] = 19;
        weight_rom[10663] = 39;
        weight_rom[10664] = 35;
        weight_rom[10665] = 19;
        weight_rom[10666] = 17;
        weight_rom[10667] = -6;
        weight_rom[10668] = 1;
        weight_rom[10669] = 2;
        weight_rom[10670] = 28;
        weight_rom[10671] = 40;
        weight_rom[10672] = 24;
        weight_rom[10673] = 30;
        weight_rom[10674] = 25;
        weight_rom[10675] = 28;
        weight_rom[10676] = 22;
        weight_rom[10677] = 14;
        weight_rom[10678] = 4;
        weight_rom[10679] = -1;
        weight_rom[10680] = 3;
        weight_rom[10681] = -8;
        weight_rom[10682] = -12;
        weight_rom[10683] = 3;
        weight_rom[10684] = 20;
        weight_rom[10685] = 26;
        weight_rom[10686] = 14;
        weight_rom[10687] = 21;
        weight_rom[10688] = 8;
        weight_rom[10689] = 14;
        weight_rom[10690] = 17;
        weight_rom[10691] = 17;
        weight_rom[10692] = 2;
        weight_rom[10693] = -4;
        weight_rom[10694] = 13;
        weight_rom[10695] = 1;
        weight_rom[10696] = 4;
        weight_rom[10697] = 3;
        weight_rom[10698] = 24;
        weight_rom[10699] = 46;
        weight_rom[10700] = 24;
        weight_rom[10701] = 43;
        weight_rom[10702] = 58;
        weight_rom[10703] = 41;
        weight_rom[10704] = 32;
        weight_rom[10705] = 15;
        weight_rom[10706] = 15;
        weight_rom[10707] = 5;
        weight_rom[10708] = 12;
        weight_rom[10709] = 4;
        weight_rom[10710] = 0;
        weight_rom[10711] = 17;
        weight_rom[10712] = 30;
        weight_rom[10713] = 24;
        weight_rom[10714] = 3;
        weight_rom[10715] = 16;
        weight_rom[10716] = 11;
        weight_rom[10717] = 15;
        weight_rom[10718] = 42;
        weight_rom[10719] = 32;
        weight_rom[10720] = 31;
        weight_rom[10721] = 7;
        weight_rom[10722] = -11;
        weight_rom[10723] = -5;
        weight_rom[10724] = 2;
        weight_rom[10725] = 7;
        weight_rom[10726] = 7;
        weight_rom[10727] = 31;
        weight_rom[10728] = 34;
        weight_rom[10729] = 74;
        weight_rom[10730] = 44;
        weight_rom[10731] = 34;
        weight_rom[10732] = 33;
        weight_rom[10733] = 24;
        weight_rom[10734] = 26;
        weight_rom[10735] = 14;
        weight_rom[10736] = 17;
        weight_rom[10737] = 17;
        weight_rom[10738] = 13;
        weight_rom[10739] = 24;
        weight_rom[10740] = 22;
        weight_rom[10741] = 21;
        weight_rom[10742] = 24;
        weight_rom[10743] = 6;
        weight_rom[10744] = 7;
        weight_rom[10745] = 26;
        weight_rom[10746] = 25;
        weight_rom[10747] = 30;
        weight_rom[10748] = -13;
        weight_rom[10749] = -14;
        weight_rom[10750] = -4;
        weight_rom[10751] = -2;
        weight_rom[10752] = 3;
        weight_rom[10753] = 15;
        weight_rom[10754] = 1;
        weight_rom[10755] = 30;
        weight_rom[10756] = 30;
        weight_rom[10757] = 45;
        weight_rom[10758] = 31;
        weight_rom[10759] = 33;
        weight_rom[10760] = 26;
        weight_rom[10761] = 25;
        weight_rom[10762] = 20;
        weight_rom[10763] = 11;
        weight_rom[10764] = 13;
        weight_rom[10765] = 16;
        weight_rom[10766] = 8;
        weight_rom[10767] = 21;
        weight_rom[10768] = 14;
        weight_rom[10769] = 12;
        weight_rom[10770] = 13;
        weight_rom[10771] = -4;
        weight_rom[10772] = 13;
        weight_rom[10773] = 21;
        weight_rom[10774] = 14;
        weight_rom[10775] = 12;
        weight_rom[10776] = -28;
        weight_rom[10777] = -7;
        weight_rom[10778] = -7;
        weight_rom[10779] = 1;
        weight_rom[10780] = 0;
        weight_rom[10781] = 2;
        weight_rom[10782] = 23;
        weight_rom[10783] = 23;
        weight_rom[10784] = 9;
        weight_rom[10785] = 7;
        weight_rom[10786] = 16;
        weight_rom[10787] = 14;
        weight_rom[10788] = 13;
        weight_rom[10789] = 14;
        weight_rom[10790] = 1;
        weight_rom[10791] = 14;
        weight_rom[10792] = 14;
        weight_rom[10793] = 26;
        weight_rom[10794] = 15;
        weight_rom[10795] = 13;
        weight_rom[10796] = 0;
        weight_rom[10797] = 7;
        weight_rom[10798] = 9;
        weight_rom[10799] = -2;
        weight_rom[10800] = -3;
        weight_rom[10801] = -8;
        weight_rom[10802] = 23;
        weight_rom[10803] = 18;
        weight_rom[10804] = -37;
        weight_rom[10805] = -18;
        weight_rom[10806] = -11;
        weight_rom[10807] = -4;
        weight_rom[10808] = -1;
        weight_rom[10809] = -2;
        weight_rom[10810] = 21;
        weight_rom[10811] = 33;
        weight_rom[10812] = 0;
        weight_rom[10813] = -29;
        weight_rom[10814] = -8;
        weight_rom[10815] = 3;
        weight_rom[10816] = -7;
        weight_rom[10817] = 2;
        weight_rom[10818] = 6;
        weight_rom[10819] = 25;
        weight_rom[10820] = 23;
        weight_rom[10821] = 30;
        weight_rom[10822] = 8;
        weight_rom[10823] = 19;
        weight_rom[10824] = 7;
        weight_rom[10825] = 6;
        weight_rom[10826] = 10;
        weight_rom[10827] = -2;
        weight_rom[10828] = 0;
        weight_rom[10829] = 10;
        weight_rom[10830] = 1;
        weight_rom[10831] = -9;
        weight_rom[10832] = -29;
        weight_rom[10833] = -10;
        weight_rom[10834] = -9;
        weight_rom[10835] = -3;
        weight_rom[10836] = 1;
        weight_rom[10837] = 1;
        weight_rom[10838] = 6;
        weight_rom[10839] = 37;
        weight_rom[10840] = 1;
        weight_rom[10841] = -16;
        weight_rom[10842] = -25;
        weight_rom[10843] = -14;
        weight_rom[10844] = 5;
        weight_rom[10845] = 19;
        weight_rom[10846] = 12;
        weight_rom[10847] = 20;
        weight_rom[10848] = 19;
        weight_rom[10849] = 20;
        weight_rom[10850] = 18;
        weight_rom[10851] = 11;
        weight_rom[10852] = 17;
        weight_rom[10853] = 8;
        weight_rom[10854] = 13;
        weight_rom[10855] = 17;
        weight_rom[10856] = 20;
        weight_rom[10857] = 3;
        weight_rom[10858] = -12;
        weight_rom[10859] = 7;
        weight_rom[10860] = -16;
        weight_rom[10861] = 21;
        weight_rom[10862] = -12;
        weight_rom[10863] = 3;
        weight_rom[10864] = 0;
        weight_rom[10865] = -1;
        weight_rom[10866] = 9;
        weight_rom[10867] = 15;
        weight_rom[10868] = 6;
        weight_rom[10869] = -36;
        weight_rom[10870] = -18;
        weight_rom[10871] = -5;
        weight_rom[10872] = -6;
        weight_rom[10873] = 17;
        weight_rom[10874] = 5;
        weight_rom[10875] = 20;
        weight_rom[10876] = 18;
        weight_rom[10877] = 19;
        weight_rom[10878] = 22;
        weight_rom[10879] = 11;
        weight_rom[10880] = 24;
        weight_rom[10881] = -2;
        weight_rom[10882] = 5;
        weight_rom[10883] = 3;
        weight_rom[10884] = -6;
        weight_rom[10885] = -1;
        weight_rom[10886] = -6;
        weight_rom[10887] = -11;
        weight_rom[10888] = 1;
        weight_rom[10889] = 20;
        weight_rom[10890] = -4;
        weight_rom[10891] = -2;
        weight_rom[10892] = 4;
        weight_rom[10893] = 2;
        weight_rom[10894] = -4;
        weight_rom[10895] = -1;
        weight_rom[10896] = -8;
        weight_rom[10897] = -27;
        weight_rom[10898] = 0;
        weight_rom[10899] = -16;
        weight_rom[10900] = -19;
        weight_rom[10901] = -19;
        weight_rom[10902] = 12;
        weight_rom[10903] = -7;
        weight_rom[10904] = -4;
        weight_rom[10905] = -2;
        weight_rom[10906] = -4;
        weight_rom[10907] = 0;
        weight_rom[10908] = -5;
        weight_rom[10909] = -11;
        weight_rom[10910] = -25;
        weight_rom[10911] = -18;
        weight_rom[10912] = -25;
        weight_rom[10913] = -27;
        weight_rom[10914] = -1;
        weight_rom[10915] = 3;
        weight_rom[10916] = 0;
        weight_rom[10917] = 1;
        weight_rom[10918] = 0;
        weight_rom[10919] = -4;
        weight_rom[10920] = 2;
        weight_rom[10921] = -1;
        weight_rom[10922] = 1;
        weight_rom[10923] = -4;
        weight_rom[10924] = -23;
        weight_rom[10925] = -14;
        weight_rom[10926] = -16;
        weight_rom[10927] = -39;
        weight_rom[10928] = -47;
        weight_rom[10929] = -40;
        weight_rom[10930] = -41;
        weight_rom[10931] = -38;
        weight_rom[10932] = -29;
        weight_rom[10933] = -44;
        weight_rom[10934] = -70;
        weight_rom[10935] = -50;
        weight_rom[10936] = -44;
        weight_rom[10937] = -32;
        weight_rom[10938] = -26;
        weight_rom[10939] = -32;
        weight_rom[10940] = -19;
        weight_rom[10941] = -20;
        weight_rom[10942] = -14;
        weight_rom[10943] = -5;
        weight_rom[10944] = -3;
        weight_rom[10945] = 3;
        weight_rom[10946] = 2;
        weight_rom[10947] = 1;
        weight_rom[10948] = 0;
        weight_rom[10949] = 3;
        weight_rom[10950] = 4;
        weight_rom[10951] = 1;
        weight_rom[10952] = -4;
        weight_rom[10953] = -15;
        weight_rom[10954] = -24;
        weight_rom[10955] = -28;
        weight_rom[10956] = -26;
        weight_rom[10957] = -23;
        weight_rom[10958] = -33;
        weight_rom[10959] = -11;
        weight_rom[10960] = -27;
        weight_rom[10961] = -36;
        weight_rom[10962] = -34;
        weight_rom[10963] = -21;
        weight_rom[10964] = -22;
        weight_rom[10965] = -13;
        weight_rom[10966] = -37;
        weight_rom[10967] = -15;
        weight_rom[10968] = -24;
        weight_rom[10969] = -19;
        weight_rom[10970] = -9;
        weight_rom[10971] = 0;
        weight_rom[10972] = -3;
        weight_rom[10973] = 0;
        weight_rom[10974] = 3;
        weight_rom[10975] = -2;
        weight_rom[10976] = -1;
        weight_rom[10977] = 2;
        weight_rom[10978] = 3;
        weight_rom[10979] = 3;
        weight_rom[10980] = -4;
        weight_rom[10981] = -1;
        weight_rom[10982] = 1;
        weight_rom[10983] = 1;
        weight_rom[10984] = 2;
        weight_rom[10985] = 4;
        weight_rom[10986] = -4;
        weight_rom[10987] = 0;
        weight_rom[10988] = -3;
        weight_rom[10989] = -4;
        weight_rom[10990] = -3;
        weight_rom[10991] = -2;
        weight_rom[10992] = 4;
        weight_rom[10993] = 3;
        weight_rom[10994] = 4;
        weight_rom[10995] = 2;
        weight_rom[10996] = -3;
        weight_rom[10997] = 3;
        weight_rom[10998] = -2;
        weight_rom[10999] = -4;
        weight_rom[11000] = 4;
        weight_rom[11001] = 1;
        weight_rom[11002] = -4;
        weight_rom[11003] = 4;
        weight_rom[11004] = -4;
        weight_rom[11005] = -2;
        weight_rom[11006] = -1;
        weight_rom[11007] = 1;
        weight_rom[11008] = 1;
        weight_rom[11009] = -3;
        weight_rom[11010] = -6;
        weight_rom[11011] = -8;
        weight_rom[11012] = -13;
        weight_rom[11013] = -10;
        weight_rom[11014] = -15;
        weight_rom[11015] = -15;
        weight_rom[11016] = -13;
        weight_rom[11017] = -19;
        weight_rom[11018] = -29;
        weight_rom[11019] = -6;
        weight_rom[11020] = -21;
        weight_rom[11021] = -28;
        weight_rom[11022] = -27;
        weight_rom[11023] = -13;
        weight_rom[11024] = -15;
        weight_rom[11025] = -10;
        weight_rom[11026] = -8;
        weight_rom[11027] = 4;
        weight_rom[11028] = 2;
        weight_rom[11029] = -3;
        weight_rom[11030] = 1;
        weight_rom[11031] = 4;
        weight_rom[11032] = -1;
        weight_rom[11033] = -2;
        weight_rom[11034] = 4;
        weight_rom[11035] = -2;
        weight_rom[11036] = -10;
        weight_rom[11037] = 0;
        weight_rom[11038] = -8;
        weight_rom[11039] = -18;
        weight_rom[11040] = -22;
        weight_rom[11041] = -7;
        weight_rom[11042] = -20;
        weight_rom[11043] = -5;
        weight_rom[11044] = -12;
        weight_rom[11045] = -5;
        weight_rom[11046] = -18;
        weight_rom[11047] = -1;
        weight_rom[11048] = -13;
        weight_rom[11049] = -23;
        weight_rom[11050] = -25;
        weight_rom[11051] = -19;
        weight_rom[11052] = -3;
        weight_rom[11053] = 4;
        weight_rom[11054] = 10;
        weight_rom[11055] = 15;
        weight_rom[11056] = 9;
        weight_rom[11057] = 13;
        weight_rom[11058] = -4;
        weight_rom[11059] = 0;
        weight_rom[11060] = 4;
        weight_rom[11061] = 1;
        weight_rom[11062] = -12;
        weight_rom[11063] = 3;
        weight_rom[11064] = -4;
        weight_rom[11065] = 20;
        weight_rom[11066] = 0;
        weight_rom[11067] = 8;
        weight_rom[11068] = 15;
        weight_rom[11069] = 0;
        weight_rom[11070] = 16;
        weight_rom[11071] = 29;
        weight_rom[11072] = 22;
        weight_rom[11073] = 3;
        weight_rom[11074] = 3;
        weight_rom[11075] = -12;
        weight_rom[11076] = -8;
        weight_rom[11077] = -23;
        weight_rom[11078] = -38;
        weight_rom[11079] = 3;
        weight_rom[11080] = -2;
        weight_rom[11081] = 3;
        weight_rom[11082] = 19;
        weight_rom[11083] = 30;
        weight_rom[11084] = 19;
        weight_rom[11085] = 9;
        weight_rom[11086] = 3;
        weight_rom[11087] = 1;
        weight_rom[11088] = 4;
        weight_rom[11089] = -2;
        weight_rom[11090] = 13;
        weight_rom[11091] = 0;
        weight_rom[11092] = 14;
        weight_rom[11093] = 27;
        weight_rom[11094] = 19;
        weight_rom[11095] = 6;
        weight_rom[11096] = 13;
        weight_rom[11097] = -5;
        weight_rom[11098] = 2;
        weight_rom[11099] = 0;
        weight_rom[11100] = 5;
        weight_rom[11101] = 11;
        weight_rom[11102] = -5;
        weight_rom[11103] = -19;
        weight_rom[11104] = -22;
        weight_rom[11105] = -30;
        weight_rom[11106] = -37;
        weight_rom[11107] = -39;
        weight_rom[11108] = -16;
        weight_rom[11109] = -23;
        weight_rom[11110] = 0;
        weight_rom[11111] = -3;
        weight_rom[11112] = -7;
        weight_rom[11113] = 10;
        weight_rom[11114] = -8;
        weight_rom[11115] = -1;
        weight_rom[11116] = -4;
        weight_rom[11117] = 1;
        weight_rom[11118] = 2;
        weight_rom[11119] = 10;
        weight_rom[11120] = 29;
        weight_rom[11121] = 21;
        weight_rom[11122] = 5;
        weight_rom[11123] = 9;
        weight_rom[11124] = 9;
        weight_rom[11125] = 16;
        weight_rom[11126] = 15;
        weight_rom[11127] = 4;
        weight_rom[11128] = 12;
        weight_rom[11129] = 7;
        weight_rom[11130] = 1;
        weight_rom[11131] = 19;
        weight_rom[11132] = -2;
        weight_rom[11133] = -24;
        weight_rom[11134] = -28;
        weight_rom[11135] = -53;
        weight_rom[11136] = -61;
        weight_rom[11137] = -27;
        weight_rom[11138] = -17;
        weight_rom[11139] = -21;
        weight_rom[11140] = -13;
        weight_rom[11141] = 8;
        weight_rom[11142] = -3;
        weight_rom[11143] = 1;
        weight_rom[11144] = 0;
        weight_rom[11145] = -1;
        weight_rom[11146] = 10;
        weight_rom[11147] = 17;
        weight_rom[11148] = 28;
        weight_rom[11149] = 5;
        weight_rom[11150] = 5;
        weight_rom[11151] = 2;
        weight_rom[11152] = 3;
        weight_rom[11153] = 13;
        weight_rom[11154] = 9;
        weight_rom[11155] = 3;
        weight_rom[11156] = -7;
        weight_rom[11157] = -3;
        weight_rom[11158] = 6;
        weight_rom[11159] = 12;
        weight_rom[11160] = 1;
        weight_rom[11161] = -14;
        weight_rom[11162] = -25;
        weight_rom[11163] = -65;
        weight_rom[11164] = -57;
        weight_rom[11165] = -28;
        weight_rom[11166] = -40;
        weight_rom[11167] = -23;
        weight_rom[11168] = -11;
        weight_rom[11169] = -16;
        weight_rom[11170] = -11;
        weight_rom[11171] = 3;
        weight_rom[11172] = 3;
        weight_rom[11173] = -1;
        weight_rom[11174] = -9;
        weight_rom[11175] = 25;
        weight_rom[11176] = 18;
        weight_rom[11177] = 3;
        weight_rom[11178] = 1;
        weight_rom[11179] = 0;
        weight_rom[11180] = -12;
        weight_rom[11181] = -14;
        weight_rom[11182] = -12;
        weight_rom[11183] = -12;
        weight_rom[11184] = -8;
        weight_rom[11185] = 8;
        weight_rom[11186] = 10;
        weight_rom[11187] = 22;
        weight_rom[11188] = 9;
        weight_rom[11189] = 9;
        weight_rom[11190] = -37;
        weight_rom[11191] = -64;
        weight_rom[11192] = -79;
        weight_rom[11193] = -71;
        weight_rom[11194] = -59;
        weight_rom[11195] = -46;
        weight_rom[11196] = -40;
        weight_rom[11197] = -21;
        weight_rom[11198] = 6;
        weight_rom[11199] = 10;
        weight_rom[11200] = -1;
        weight_rom[11201] = 0;
        weight_rom[11202] = 22;
        weight_rom[11203] = 10;
        weight_rom[11204] = 20;
        weight_rom[11205] = -7;
        weight_rom[11206] = -7;
        weight_rom[11207] = -7;
        weight_rom[11208] = -15;
        weight_rom[11209] = -14;
        weight_rom[11210] = 6;
        weight_rom[11211] = -15;
        weight_rom[11212] = -3;
        weight_rom[11213] = 19;
        weight_rom[11214] = 31;
        weight_rom[11215] = 49;
        weight_rom[11216] = 32;
        weight_rom[11217] = 13;
        weight_rom[11218] = -39;
        weight_rom[11219] = -60;
        weight_rom[11220] = -72;
        weight_rom[11221] = -67;
        weight_rom[11222] = -57;
        weight_rom[11223] = -50;
        weight_rom[11224] = -36;
        weight_rom[11225] = -34;
        weight_rom[11226] = 2;
        weight_rom[11227] = 4;
        weight_rom[11228] = 13;
        weight_rom[11229] = 16;
        weight_rom[11230] = 34;
        weight_rom[11231] = 14;
        weight_rom[11232] = 13;
        weight_rom[11233] = -6;
        weight_rom[11234] = -13;
        weight_rom[11235] = -7;
        weight_rom[11236] = -24;
        weight_rom[11237] = -7;
        weight_rom[11238] = -22;
        weight_rom[11239] = -12;
        weight_rom[11240] = 3;
        weight_rom[11241] = 34;
        weight_rom[11242] = 67;
        weight_rom[11243] = 68;
        weight_rom[11244] = 34;
        weight_rom[11245] = 6;
        weight_rom[11246] = -43;
        weight_rom[11247] = -53;
        weight_rom[11248] = -70;
        weight_rom[11249] = -64;
        weight_rom[11250] = -52;
        weight_rom[11251] = -45;
        weight_rom[11252] = -29;
        weight_rom[11253] = -24;
        weight_rom[11254] = 4;
        weight_rom[11255] = 7;
        weight_rom[11256] = 14;
        weight_rom[11257] = 13;
        weight_rom[11258] = 28;
        weight_rom[11259] = 9;
        weight_rom[11260] = 7;
        weight_rom[11261] = -1;
        weight_rom[11262] = -6;
        weight_rom[11263] = -7;
        weight_rom[11264] = -22;
        weight_rom[11265] = -24;
        weight_rom[11266] = -17;
        weight_rom[11267] = 4;
        weight_rom[11268] = 17;
        weight_rom[11269] = 51;
        weight_rom[11270] = 71;
        weight_rom[11271] = 52;
        weight_rom[11272] = 35;
        weight_rom[11273] = -12;
        weight_rom[11274] = -51;
        weight_rom[11275] = -60;
        weight_rom[11276] = -64;
        weight_rom[11277] = -49;
        weight_rom[11278] = -27;
        weight_rom[11279] = -38;
        weight_rom[11280] = -36;
        weight_rom[11281] = -13;
        weight_rom[11282] = 3;
        weight_rom[11283] = -5;
        weight_rom[11284] = 2;
        weight_rom[11285] = 20;
        weight_rom[11286] = 26;
        weight_rom[11287] = 18;
        weight_rom[11288] = -5;
        weight_rom[11289] = -8;
        weight_rom[11290] = -11;
        weight_rom[11291] = -12;
        weight_rom[11292] = -21;
        weight_rom[11293] = 2;
        weight_rom[11294] = 11;
        weight_rom[11295] = 13;
        weight_rom[11296] = 23;
        weight_rom[11297] = 48;
        weight_rom[11298] = 56;
        weight_rom[11299] = 29;
        weight_rom[11300] = -2;
        weight_rom[11301] = -42;
        weight_rom[11302] = -63;
        weight_rom[11303] = -52;
        weight_rom[11304] = -33;
        weight_rom[11305] = -25;
        weight_rom[11306] = -23;
        weight_rom[11307] = -20;
        weight_rom[11308] = -29;
        weight_rom[11309] = -7;
        weight_rom[11310] = -18;
        weight_rom[11311] = -8;
        weight_rom[11312] = -1;
        weight_rom[11313] = -1;
        weight_rom[11314] = 15;
        weight_rom[11315] = 3;
        weight_rom[11316] = -11;
        weight_rom[11317] = 0;
        weight_rom[11318] = -19;
        weight_rom[11319] = -3;
        weight_rom[11320] = 0;
        weight_rom[11321] = 9;
        weight_rom[11322] = 1;
        weight_rom[11323] = 2;
        weight_rom[11324] = 33;
        weight_rom[11325] = 38;
        weight_rom[11326] = 42;
        weight_rom[11327] = 13;
        weight_rom[11328] = -9;
        weight_rom[11329] = -35;
        weight_rom[11330] = -27;
        weight_rom[11331] = -25;
        weight_rom[11332] = -22;
        weight_rom[11333] = -3;
        weight_rom[11334] = -8;
        weight_rom[11335] = -6;
        weight_rom[11336] = 9;
        weight_rom[11337] = 17;
        weight_rom[11338] = -15;
        weight_rom[11339] = -9;
        weight_rom[11340] = 0;
        weight_rom[11341] = 4;
        weight_rom[11342] = 5;
        weight_rom[11343] = 0;
        weight_rom[11344] = -4;
        weight_rom[11345] = -18;
        weight_rom[11346] = -4;
        weight_rom[11347] = 0;
        weight_rom[11348] = 0;
        weight_rom[11349] = 9;
        weight_rom[11350] = 2;
        weight_rom[11351] = 5;
        weight_rom[11352] = 15;
        weight_rom[11353] = 19;
        weight_rom[11354] = 20;
        weight_rom[11355] = 1;
        weight_rom[11356] = -8;
        weight_rom[11357] = -18;
        weight_rom[11358] = -20;
        weight_rom[11359] = -13;
        weight_rom[11360] = -9;
        weight_rom[11361] = -5;
        weight_rom[11362] = -8;
        weight_rom[11363] = 14;
        weight_rom[11364] = 24;
        weight_rom[11365] = 32;
        weight_rom[11366] = 20;
        weight_rom[11367] = 10;
        weight_rom[11368] = -1;
        weight_rom[11369] = 9;
        weight_rom[11370] = 17;
        weight_rom[11371] = 6;
        weight_rom[11372] = -3;
        weight_rom[11373] = -8;
        weight_rom[11374] = -10;
        weight_rom[11375] = -23;
        weight_rom[11376] = -2;
        weight_rom[11377] = 13;
        weight_rom[11378] = -13;
        weight_rom[11379] = -9;
        weight_rom[11380] = 13;
        weight_rom[11381] = 10;
        weight_rom[11382] = 21;
        weight_rom[11383] = 5;
        weight_rom[11384] = -4;
        weight_rom[11385] = -9;
        weight_rom[11386] = -4;
        weight_rom[11387] = -4;
        weight_rom[11388] = -11;
        weight_rom[11389] = 1;
        weight_rom[11390] = -3;
        weight_rom[11391] = 21;
        weight_rom[11392] = 5;
        weight_rom[11393] = 9;
        weight_rom[11394] = 16;
        weight_rom[11395] = -1;
        weight_rom[11396] = -4;
        weight_rom[11397] = 1;
        weight_rom[11398] = -4;
        weight_rom[11399] = 12;
        weight_rom[11400] = -1;
        weight_rom[11401] = 9;
        weight_rom[11402] = -16;
        weight_rom[11403] = -19;
        weight_rom[11404] = -5;
        weight_rom[11405] = 5;
        weight_rom[11406] = -1;
        weight_rom[11407] = 8;
        weight_rom[11408] = 4;
        weight_rom[11409] = 8;
        weight_rom[11410] = 15;
        weight_rom[11411] = 7;
        weight_rom[11412] = -1;
        weight_rom[11413] = -6;
        weight_rom[11414] = -9;
        weight_rom[11415] = -5;
        weight_rom[11416] = 4;
        weight_rom[11417] = 12;
        weight_rom[11418] = 17;
        weight_rom[11419] = 14;
        weight_rom[11420] = 3;
        weight_rom[11421] = -13;
        weight_rom[11422] = 26;
        weight_rom[11423] = 10;
        weight_rom[11424] = -2;
        weight_rom[11425] = 0;
        weight_rom[11426] = 5;
        weight_rom[11427] = 8;
        weight_rom[11428] = -3;
        weight_rom[11429] = -8;
        weight_rom[11430] = -5;
        weight_rom[11431] = 8;
        weight_rom[11432] = -4;
        weight_rom[11433] = 17;
        weight_rom[11434] = 14;
        weight_rom[11435] = 10;
        weight_rom[11436] = 0;
        weight_rom[11437] = 9;
        weight_rom[11438] = 12;
        weight_rom[11439] = -7;
        weight_rom[11440] = -3;
        weight_rom[11441] = -21;
        weight_rom[11442] = 4;
        weight_rom[11443] = -1;
        weight_rom[11444] = 8;
        weight_rom[11445] = 6;
        weight_rom[11446] = -1;
        weight_rom[11447] = 10;
        weight_rom[11448] = 9;
        weight_rom[11449] = -6;
        weight_rom[11450] = 16;
        weight_rom[11451] = 5;
        weight_rom[11452] = -1;
        weight_rom[11453] = 4;
        weight_rom[11454] = -3;
        weight_rom[11455] = 5;
        weight_rom[11456] = -10;
        weight_rom[11457] = -19;
        weight_rom[11458] = -6;
        weight_rom[11459] = -3;
        weight_rom[11460] = 2;
        weight_rom[11461] = 8;
        weight_rom[11462] = 1;
        weight_rom[11463] = -9;
        weight_rom[11464] = 0;
        weight_rom[11465] = 3;
        weight_rom[11466] = 19;
        weight_rom[11467] = -1;
        weight_rom[11468] = -4;
        weight_rom[11469] = -14;
        weight_rom[11470] = -5;
        weight_rom[11471] = 5;
        weight_rom[11472] = 11;
        weight_rom[11473] = 22;
        weight_rom[11474] = 14;
        weight_rom[11475] = 11;
        weight_rom[11476] = -4;
        weight_rom[11477] = 12;
        weight_rom[11478] = 3;
        weight_rom[11479] = 4;
        weight_rom[11480] = 4;
        weight_rom[11481] = -1;
        weight_rom[11482] = 7;
        weight_rom[11483] = 9;
        weight_rom[11484] = -12;
        weight_rom[11485] = -18;
        weight_rom[11486] = -13;
        weight_rom[11487] = -6;
        weight_rom[11488] = -6;
        weight_rom[11489] = -1;
        weight_rom[11490] = -4;
        weight_rom[11491] = -6;
        weight_rom[11492] = -1;
        weight_rom[11493] = 0;
        weight_rom[11494] = -4;
        weight_rom[11495] = 8;
        weight_rom[11496] = -1;
        weight_rom[11497] = -2;
        weight_rom[11498] = -9;
        weight_rom[11499] = 7;
        weight_rom[11500] = 10;
        weight_rom[11501] = 10;
        weight_rom[11502] = 12;
        weight_rom[11503] = 8;
        weight_rom[11504] = 4;
        weight_rom[11505] = 10;
        weight_rom[11506] = 18;
        weight_rom[11507] = 8;
        weight_rom[11508] = -2;
        weight_rom[11509] = 1;
        weight_rom[11510] = -10;
        weight_rom[11511] = 0;
        weight_rom[11512] = -7;
        weight_rom[11513] = 9;
        weight_rom[11514] = -4;
        weight_rom[11515] = -7;
        weight_rom[11516] = -10;
        weight_rom[11517] = -11;
        weight_rom[11518] = -7;
        weight_rom[11519] = -9;
        weight_rom[11520] = -13;
        weight_rom[11521] = -2;
        weight_rom[11522] = 9;
        weight_rom[11523] = -1;
        weight_rom[11524] = 4;
        weight_rom[11525] = 0;
        weight_rom[11526] = 24;
        weight_rom[11527] = 14;
        weight_rom[11528] = 7;
        weight_rom[11529] = 11;
        weight_rom[11530] = 5;
        weight_rom[11531] = 12;
        weight_rom[11532] = 1;
        weight_rom[11533] = 23;
        weight_rom[11534] = 20;
        weight_rom[11535] = 7;
        weight_rom[11536] = -3;
        weight_rom[11537] = 3;
        weight_rom[11538] = 1;
        weight_rom[11539] = -11;
        weight_rom[11540] = -24;
        weight_rom[11541] = -9;
        weight_rom[11542] = 0;
        weight_rom[11543] = 13;
        weight_rom[11544] = -7;
        weight_rom[11545] = 7;
        weight_rom[11546] = -7;
        weight_rom[11547] = -9;
        weight_rom[11548] = -3;
        weight_rom[11549] = -1;
        weight_rom[11550] = 13;
        weight_rom[11551] = 7;
        weight_rom[11552] = 5;
        weight_rom[11553] = 6;
        weight_rom[11554] = 14;
        weight_rom[11555] = 9;
        weight_rom[11556] = -1;
        weight_rom[11557] = -5;
        weight_rom[11558] = -2;
        weight_rom[11559] = -9;
        weight_rom[11560] = 11;
        weight_rom[11561] = 4;
        weight_rom[11562] = 4;
        weight_rom[11563] = 0;
        weight_rom[11564] = 3;
        weight_rom[11565] = 1;
        weight_rom[11566] = 13;
        weight_rom[11567] = 1;
        weight_rom[11568] = -11;
        weight_rom[11569] = -31;
        weight_rom[11570] = -15;
        weight_rom[11571] = -10;
        weight_rom[11572] = -14;
        weight_rom[11573] = -11;
        weight_rom[11574] = -18;
        weight_rom[11575] = -4;
        weight_rom[11576] = -12;
        weight_rom[11577] = -6;
        weight_rom[11578] = -2;
        weight_rom[11579] = 5;
        weight_rom[11580] = 6;
        weight_rom[11581] = -9;
        weight_rom[11582] = 5;
        weight_rom[11583] = 1;
        weight_rom[11584] = -13;
        weight_rom[11585] = -7;
        weight_rom[11586] = -1;
        weight_rom[11587] = -10;
        weight_rom[11588] = -6;
        weight_rom[11589] = 10;
        weight_rom[11590] = -6;
        weight_rom[11591] = 4;
        weight_rom[11592] = 2;
        weight_rom[11593] = -2;
        weight_rom[11594] = 15;
        weight_rom[11595] = 30;
        weight_rom[11596] = 11;
        weight_rom[11597] = -13;
        weight_rom[11598] = -9;
        weight_rom[11599] = -13;
        weight_rom[11600] = -7;
        weight_rom[11601] = -8;
        weight_rom[11602] = -6;
        weight_rom[11603] = -8;
        weight_rom[11604] = -23;
        weight_rom[11605] = -3;
        weight_rom[11606] = -3;
        weight_rom[11607] = -7;
        weight_rom[11608] = 1;
        weight_rom[11609] = -7;
        weight_rom[11610] = 7;
        weight_rom[11611] = 6;
        weight_rom[11612] = 6;
        weight_rom[11613] = -10;
        weight_rom[11614] = -11;
        weight_rom[11615] = -14;
        weight_rom[11616] = -6;
        weight_rom[11617] = -4;
        weight_rom[11618] = 8;
        weight_rom[11619] = -1;
        weight_rom[11620] = 2;
        weight_rom[11621] = 3;
        weight_rom[11622] = 11;
        weight_rom[11623] = 10;
        weight_rom[11624] = 15;
        weight_rom[11625] = -11;
        weight_rom[11626] = -11;
        weight_rom[11627] = 1;
        weight_rom[11628] = -7;
        weight_rom[11629] = -7;
        weight_rom[11630] = -9;
        weight_rom[11631] = -6;
        weight_rom[11632] = -2;
        weight_rom[11633] = 1;
        weight_rom[11634] = -6;
        weight_rom[11635] = 0;
        weight_rom[11636] = -1;
        weight_rom[11637] = 12;
        weight_rom[11638] = 7;
        weight_rom[11639] = 0;
        weight_rom[11640] = 1;
        weight_rom[11641] = -10;
        weight_rom[11642] = -20;
        weight_rom[11643] = -14;
        weight_rom[11644] = 1;
        weight_rom[11645] = -1;
        weight_rom[11646] = 11;
        weight_rom[11647] = -1;
        weight_rom[11648] = -1;
        weight_rom[11649] = -4;
        weight_rom[11650] = -4;
        weight_rom[11651] = 14;
        weight_rom[11652] = 7;
        weight_rom[11653] = 26;
        weight_rom[11654] = -7;
        weight_rom[11655] = 2;
        weight_rom[11656] = -6;
        weight_rom[11657] = 1;
        weight_rom[11658] = -1;
        weight_rom[11659] = -14;
        weight_rom[11660] = -6;
        weight_rom[11661] = 3;
        weight_rom[11662] = 5;
        weight_rom[11663] = -11;
        weight_rom[11664] = 8;
        weight_rom[11665] = 13;
        weight_rom[11666] = 11;
        weight_rom[11667] = 2;
        weight_rom[11668] = -2;
        weight_rom[11669] = -12;
        weight_rom[11670] = -11;
        weight_rom[11671] = -17;
        weight_rom[11672] = 2;
        weight_rom[11673] = 10;
        weight_rom[11674] = 4;
        weight_rom[11675] = -1;
        weight_rom[11676] = 3;
        weight_rom[11677] = -4;
        weight_rom[11678] = 2;
        weight_rom[11679] = 2;
        weight_rom[11680] = 5;
        weight_rom[11681] = 8;
        weight_rom[11682] = 28;
        weight_rom[11683] = 14;
        weight_rom[11684] = 10;
        weight_rom[11685] = -12;
        weight_rom[11686] = -16;
        weight_rom[11687] = -10;
        weight_rom[11688] = -15;
        weight_rom[11689] = 4;
        weight_rom[11690] = 4;
        weight_rom[11691] = -13;
        weight_rom[11692] = -16;
        weight_rom[11693] = -8;
        weight_rom[11694] = -2;
        weight_rom[11695] = -1;
        weight_rom[11696] = 2;
        weight_rom[11697] = -8;
        weight_rom[11698] = -9;
        weight_rom[11699] = -19;
        weight_rom[11700] = -3;
        weight_rom[11701] = 0;
        weight_rom[11702] = 1;
        weight_rom[11703] = 1;
        weight_rom[11704] = 1;
        weight_rom[11705] = 0;
        weight_rom[11706] = 3;
        weight_rom[11707] = -4;
        weight_rom[11708] = 4;
        weight_rom[11709] = -3;
        weight_rom[11710] = 0;
        weight_rom[11711] = 1;
        weight_rom[11712] = 5;
        weight_rom[11713] = -17;
        weight_rom[11714] = -8;
        weight_rom[11715] = -10;
        weight_rom[11716] = -27;
        weight_rom[11717] = -34;
        weight_rom[11718] = -29;
        weight_rom[11719] = -16;
        weight_rom[11720] = -34;
        weight_rom[11721] = -1;
        weight_rom[11722] = 1;
        weight_rom[11723] = 16;
        weight_rom[11724] = 10;
        weight_rom[11725] = 0;
        weight_rom[11726] = -21;
        weight_rom[11727] = -6;
        weight_rom[11728] = 3;
        weight_rom[11729] = 4;
        weight_rom[11730] = 3;
        weight_rom[11731] = -1;
        weight_rom[11732] = 2;
        weight_rom[11733] = 2;
        weight_rom[11734] = -2;
        weight_rom[11735] = -2;
        weight_rom[11736] = 2;
        weight_rom[11737] = -4;
        weight_rom[11738] = -2;
        weight_rom[11739] = 1;
        weight_rom[11740] = 1;
        weight_rom[11741] = 0;
        weight_rom[11742] = 3;
        weight_rom[11743] = -7;
        weight_rom[11744] = 6;
        weight_rom[11745] = 9;
        weight_rom[11746] = -1;
        weight_rom[11747] = -8;
        weight_rom[11748] = 10;
        weight_rom[11749] = 32;
        weight_rom[11750] = 10;
        weight_rom[11751] = -5;
        weight_rom[11752] = 13;
        weight_rom[11753] = 5;
        weight_rom[11754] = -4;
        weight_rom[11755] = 1;
        weight_rom[11756] = 4;
        weight_rom[11757] = 3;
        weight_rom[11758] = 2;
        weight_rom[11759] = -3;
        weight_rom[11760] = -4;
        weight_rom[11761] = -3;
        weight_rom[11762] = 1;
        weight_rom[11763] = -4;
        weight_rom[11764] = 1;
        weight_rom[11765] = -3;
        weight_rom[11766] = 1;
        weight_rom[11767] = -1;
        weight_rom[11768] = -4;
        weight_rom[11769] = 4;
        weight_rom[11770] = 1;
        weight_rom[11771] = 1;
        weight_rom[11772] = -3;
        weight_rom[11773] = -2;
        weight_rom[11774] = 5;
        weight_rom[11775] = 2;
        weight_rom[11776] = 2;
        weight_rom[11777] = 1;
        weight_rom[11778] = 2;
        weight_rom[11779] = 1;
        weight_rom[11780] = -1;
        weight_rom[11781] = -4;
        weight_rom[11782] = 2;
        weight_rom[11783] = -4;
        weight_rom[11784] = 4;
        weight_rom[11785] = -4;
        weight_rom[11786] = -2;
        weight_rom[11787] = -1;
        weight_rom[11788] = -4;
        weight_rom[11789] = 2;
        weight_rom[11790] = 4;
        weight_rom[11791] = 3;
        weight_rom[11792] = 3;
        weight_rom[11793] = 1;
        weight_rom[11794] = 18;
        weight_rom[11795] = 20;
        weight_rom[11796] = 15;
        weight_rom[11797] = 1;
        weight_rom[11798] = 4;
        weight_rom[11799] = -5;
        weight_rom[11800] = 5;
        weight_rom[11801] = 17;
        weight_rom[11802] = 8;
        weight_rom[11803] = 19;
        weight_rom[11804] = 3;
        weight_rom[11805] = 14;
        weight_rom[11806] = 3;
        weight_rom[11807] = 23;
        weight_rom[11808] = 20;
        weight_rom[11809] = 15;
        weight_rom[11810] = 14;
        weight_rom[11811] = 14;
        weight_rom[11812] = 1;
        weight_rom[11813] = 4;
        weight_rom[11814] = 4;
        weight_rom[11815] = -3;
        weight_rom[11816] = 4;
        weight_rom[11817] = 3;
        weight_rom[11818] = 4;
        weight_rom[11819] = 2;
        weight_rom[11820] = -13;
        weight_rom[11821] = -1;
        weight_rom[11822] = 17;
        weight_rom[11823] = 25;
        weight_rom[11824] = 26;
        weight_rom[11825] = 43;
        weight_rom[11826] = 39;
        weight_rom[11827] = 45;
        weight_rom[11828] = 45;
        weight_rom[11829] = 43;
        weight_rom[11830] = 64;
        weight_rom[11831] = 49;
        weight_rom[11832] = 40;
        weight_rom[11833] = 15;
        weight_rom[11834] = 5;
        weight_rom[11835] = 6;
        weight_rom[11836] = 22;
        weight_rom[11837] = 12;
        weight_rom[11838] = 21;
        weight_rom[11839] = 24;
        weight_rom[11840] = 32;
        weight_rom[11841] = 14;
        weight_rom[11842] = 4;
        weight_rom[11843] = 2;
        weight_rom[11844] = 4;
        weight_rom[11845] = -2;
        weight_rom[11846] = 10;
        weight_rom[11847] = -4;
        weight_rom[11848] = 3;
        weight_rom[11849] = 19;
        weight_rom[11850] = 36;
        weight_rom[11851] = 35;
        weight_rom[11852] = 18;
        weight_rom[11853] = 36;
        weight_rom[11854] = 34;
        weight_rom[11855] = 27;
        weight_rom[11856] = 26;
        weight_rom[11857] = 25;
        weight_rom[11858] = 13;
        weight_rom[11859] = 25;
        weight_rom[11860] = 13;
        weight_rom[11861] = 8;
        weight_rom[11862] = 9;
        weight_rom[11863] = 11;
        weight_rom[11864] = -5;
        weight_rom[11865] = 2;
        weight_rom[11866] = -9;
        weight_rom[11867] = 7;
        weight_rom[11868] = 14;
        weight_rom[11869] = -13;
        weight_rom[11870] = 4;
        weight_rom[11871] = -3;
        weight_rom[11872] = 4;
        weight_rom[11873] = 3;
        weight_rom[11874] = 9;
        weight_rom[11875] = -4;
        weight_rom[11876] = 3;
        weight_rom[11877] = 31;
        weight_rom[11878] = 47;
        weight_rom[11879] = 26;
        weight_rom[11880] = 28;
        weight_rom[11881] = 22;
        weight_rom[11882] = 29;
        weight_rom[11883] = 7;
        weight_rom[11884] = 25;
        weight_rom[11885] = 29;
        weight_rom[11886] = 17;
        weight_rom[11887] = 5;
        weight_rom[11888] = 20;
        weight_rom[11889] = 19;
        weight_rom[11890] = 12;
        weight_rom[11891] = 10;
        weight_rom[11892] = 16;
        weight_rom[11893] = -13;
        weight_rom[11894] = -8;
        weight_rom[11895] = -15;
        weight_rom[11896] = -28;
        weight_rom[11897] = -4;
        weight_rom[11898] = -5;
        weight_rom[11899] = -1;
        weight_rom[11900] = 4;
        weight_rom[11901] = -1;
        weight_rom[11902] = 3;
        weight_rom[11903] = 9;
        weight_rom[11904] = 35;
        weight_rom[11905] = 31;
        weight_rom[11906] = 29;
        weight_rom[11907] = 31;
        weight_rom[11908] = 20;
        weight_rom[11909] = 17;
        weight_rom[11910] = 12;
        weight_rom[11911] = -1;
        weight_rom[11912] = 13;
        weight_rom[11913] = 10;
        weight_rom[11914] = 20;
        weight_rom[11915] = 11;
        weight_rom[11916] = 27;
        weight_rom[11917] = 13;
        weight_rom[11918] = 18;
        weight_rom[11919] = 17;
        weight_rom[11920] = 7;
        weight_rom[11921] = 11;
        weight_rom[11922] = 19;
        weight_rom[11923] = 14;
        weight_rom[11924] = 5;
        weight_rom[11925] = -22;
        weight_rom[11926] = 0;
        weight_rom[11927] = -2;
        weight_rom[11928] = 0;
        weight_rom[11929] = 0;
        weight_rom[11930] = -17;
        weight_rom[11931] = 15;
        weight_rom[11932] = 17;
        weight_rom[11933] = 30;
        weight_rom[11934] = 31;
        weight_rom[11935] = 24;
        weight_rom[11936] = 8;
        weight_rom[11937] = 21;
        weight_rom[11938] = 2;
        weight_rom[11939] = -2;
        weight_rom[11940] = -5;
        weight_rom[11941] = -10;
        weight_rom[11942] = -13;
        weight_rom[11943] = -10;
        weight_rom[11944] = -9;
        weight_rom[11945] = -7;
        weight_rom[11946] = -10;
        weight_rom[11947] = -4;
        weight_rom[11948] = -3;
        weight_rom[11949] = -1;
        weight_rom[11950] = 14;
        weight_rom[11951] = 23;
        weight_rom[11952] = -4;
        weight_rom[11953] = -10;
        weight_rom[11954] = -8;
        weight_rom[11955] = 14;
        weight_rom[11956] = 3;
        weight_rom[11957] = 21;
        weight_rom[11958] = 15;
        weight_rom[11959] = 25;
        weight_rom[11960] = 59;
        weight_rom[11961] = 42;
        weight_rom[11962] = 25;
        weight_rom[11963] = 18;
        weight_rom[11964] = 10;
        weight_rom[11965] = 0;
        weight_rom[11966] = 8;
        weight_rom[11967] = -16;
        weight_rom[11968] = -13;
        weight_rom[11969] = -16;
        weight_rom[11970] = -28;
        weight_rom[11971] = -33;
        weight_rom[11972] = -27;
        weight_rom[11973] = -21;
        weight_rom[11974] = 0;
        weight_rom[11975] = 2;
        weight_rom[11976] = 9;
        weight_rom[11977] = 13;
        weight_rom[11978] = 20;
        weight_rom[11979] = -3;
        weight_rom[11980] = -12;
        weight_rom[11981] = -15;
        weight_rom[11982] = 9;
        weight_rom[11983] = -1;
        weight_rom[11984] = 1;
        weight_rom[11985] = 6;
        weight_rom[11986] = 17;
        weight_rom[11987] = 38;
        weight_rom[11988] = 69;
        weight_rom[11989] = 25;
        weight_rom[11990] = 21;
        weight_rom[11991] = 28;
        weight_rom[11992] = 7;
        weight_rom[11993] = 13;
        weight_rom[11994] = 2;
        weight_rom[11995] = 2;
        weight_rom[11996] = 8;
        weight_rom[11997] = -7;
        weight_rom[11998] = -22;
        weight_rom[11999] = -20;
        weight_rom[12000] = -23;
        weight_rom[12001] = 1;
        weight_rom[12002] = 5;
        weight_rom[12003] = 9;
        weight_rom[12004] = 1;
        weight_rom[12005] = 2;
        weight_rom[12006] = 3;
        weight_rom[12007] = -12;
        weight_rom[12008] = -42;
        weight_rom[12009] = -28;
        weight_rom[12010] = -11;
        weight_rom[12011] = 4;
        weight_rom[12012] = 4;
        weight_rom[12013] = 6;
        weight_rom[12014] = 2;
        weight_rom[12015] = 16;
        weight_rom[12016] = 42;
        weight_rom[12017] = 27;
        weight_rom[12018] = 9;
        weight_rom[12019] = 11;
        weight_rom[12020] = 9;
        weight_rom[12021] = 6;
        weight_rom[12022] = 0;
        weight_rom[12023] = 2;
        weight_rom[12024] = -5;
        weight_rom[12025] = -18;
        weight_rom[12026] = -31;
        weight_rom[12027] = -31;
        weight_rom[12028] = -13;
        weight_rom[12029] = 4;
        weight_rom[12030] = 6;
        weight_rom[12031] = 6;
        weight_rom[12032] = 3;
        weight_rom[12033] = 8;
        weight_rom[12034] = -1;
        weight_rom[12035] = -10;
        weight_rom[12036] = -57;
        weight_rom[12037] = -46;
        weight_rom[12038] = -18;
        weight_rom[12039] = -14;
        weight_rom[12040] = 9;
        weight_rom[12041] = 7;
        weight_rom[12042] = -9;
        weight_rom[12043] = 22;
        weight_rom[12044] = 8;
        weight_rom[12045] = 8;
        weight_rom[12046] = -1;
        weight_rom[12047] = -3;
        weight_rom[12048] = 4;
        weight_rom[12049] = -9;
        weight_rom[12050] = -4;
        weight_rom[12051] = -16;
        weight_rom[12052] = -27;
        weight_rom[12053] = -34;
        weight_rom[12054] = -36;
        weight_rom[12055] = -13;
        weight_rom[12056] = 0;
        weight_rom[12057] = 19;
        weight_rom[12058] = 3;
        weight_rom[12059] = 14;
        weight_rom[12060] = -7;
        weight_rom[12061] = 2;
        weight_rom[12062] = 1;
        weight_rom[12063] = -44;
        weight_rom[12064] = -61;
        weight_rom[12065] = -55;
        weight_rom[12066] = -25;
        weight_rom[12067] = -4;
        weight_rom[12068] = 3;
        weight_rom[12069] = 3;
        weight_rom[12070] = 5;
        weight_rom[12071] = 4;
        weight_rom[12072] = -7;
        weight_rom[12073] = 2;
        weight_rom[12074] = -19;
        weight_rom[12075] = -3;
        weight_rom[12076] = -7;
        weight_rom[12077] = -6;
        weight_rom[12078] = -18;
        weight_rom[12079] = -24;
        weight_rom[12080] = -29;
        weight_rom[12081] = -39;
        weight_rom[12082] = -17;
        weight_rom[12083] = 1;
        weight_rom[12084] = 20;
        weight_rom[12085] = -4;
        weight_rom[12086] = 0;
        weight_rom[12087] = 12;
        weight_rom[12088] = 3;
        weight_rom[12089] = 3;
        weight_rom[12090] = 14;
        weight_rom[12091] = -3;
        weight_rom[12092] = -16;
        weight_rom[12093] = -36;
        weight_rom[12094] = -30;
        weight_rom[12095] = 17;
        weight_rom[12096] = 2;
        weight_rom[12097] = 14;
        weight_rom[12098] = 0;
        weight_rom[12099] = -11;
        weight_rom[12100] = -32;
        weight_rom[12101] = -25;
        weight_rom[12102] = -39;
        weight_rom[12103] = -9;
        weight_rom[12104] = -7;
        weight_rom[12105] = -7;
        weight_rom[12106] = -16;
        weight_rom[12107] = -16;
        weight_rom[12108] = -16;
        weight_rom[12109] = -17;
        weight_rom[12110] = 0;
        weight_rom[12111] = 11;
        weight_rom[12112] = 28;
        weight_rom[12113] = 12;
        weight_rom[12114] = 3;
        weight_rom[12115] = 9;
        weight_rom[12116] = 18;
        weight_rom[12117] = 24;
        weight_rom[12118] = 23;
        weight_rom[12119] = 17;
        weight_rom[12120] = 30;
        weight_rom[12121] = 22;
        weight_rom[12122] = -3;
        weight_rom[12123] = 13;
        weight_rom[12124] = -2;
        weight_rom[12125] = 9;
        weight_rom[12126] = -4;
        weight_rom[12127] = -29;
        weight_rom[12128] = -47;
        weight_rom[12129] = -44;
        weight_rom[12130] = -33;
        weight_rom[12131] = -39;
        weight_rom[12132] = -11;
        weight_rom[12133] = -13;
        weight_rom[12134] = -17;
        weight_rom[12135] = -10;
        weight_rom[12136] = -4;
        weight_rom[12137] = 16;
        weight_rom[12138] = 30;
        weight_rom[12139] = 39;
        weight_rom[12140] = 28;
        weight_rom[12141] = 13;
        weight_rom[12142] = -4;
        weight_rom[12143] = 5;
        weight_rom[12144] = 11;
        weight_rom[12145] = 15;
        weight_rom[12146] = 8;
        weight_rom[12147] = 21;
        weight_rom[12148] = 29;
        weight_rom[12149] = 35;
        weight_rom[12150] = 42;
        weight_rom[12151] = 22;
        weight_rom[12152] = 2;
        weight_rom[12153] = -1;
        weight_rom[12154] = 4;
        weight_rom[12155] = -26;
        weight_rom[12156] = -37;
        weight_rom[12157] = -21;
        weight_rom[12158] = -20;
        weight_rom[12159] = -19;
        weight_rom[12160] = -13;
        weight_rom[12161] = -14;
        weight_rom[12162] = -15;
        weight_rom[12163] = 9;
        weight_rom[12164] = 23;
        weight_rom[12165] = 31;
        weight_rom[12166] = 51;
        weight_rom[12167] = 40;
        weight_rom[12168] = 32;
        weight_rom[12169] = 15;
        weight_rom[12170] = 9;
        weight_rom[12171] = 9;
        weight_rom[12172] = 2;
        weight_rom[12173] = 5;
        weight_rom[12174] = -4;
        weight_rom[12175] = -2;
        weight_rom[12176] = -3;
        weight_rom[12177] = 33;
        weight_rom[12178] = 47;
        weight_rom[12179] = 3;
        weight_rom[12180] = -3;
        weight_rom[12181] = -6;
        weight_rom[12182] = 0;
        weight_rom[12183] = 0;
        weight_rom[12184] = -18;
        weight_rom[12185] = -13;
        weight_rom[12186] = -4;
        weight_rom[12187] = -18;
        weight_rom[12188] = -7;
        weight_rom[12189] = -17;
        weight_rom[12190] = -7;
        weight_rom[12191] = 13;
        weight_rom[12192] = 30;
        weight_rom[12193] = 52;
        weight_rom[12194] = 61;
        weight_rom[12195] = 43;
        weight_rom[12196] = 37;
        weight_rom[12197] = 14;
        weight_rom[12198] = -8;
        weight_rom[12199] = -1;
        weight_rom[12200] = -12;
        weight_rom[12201] = 0;
        weight_rom[12202] = 3;
        weight_rom[12203] = -15;
        weight_rom[12204] = 2;
        weight_rom[12205] = 33;
        weight_rom[12206] = 41;
        weight_rom[12207] = 19;
        weight_rom[12208] = -3;
        weight_rom[12209] = 3;
        weight_rom[12210] = -4;
        weight_rom[12211] = 7;
        weight_rom[12212] = -7;
        weight_rom[12213] = 5;
        weight_rom[12214] = 2;
        weight_rom[12215] = 4;
        weight_rom[12216] = -4;
        weight_rom[12217] = 8;
        weight_rom[12218] = 2;
        weight_rom[12219] = 9;
        weight_rom[12220] = 30;
        weight_rom[12221] = 42;
        weight_rom[12222] = 57;
        weight_rom[12223] = 44;
        weight_rom[12224] = 22;
        weight_rom[12225] = 5;
        weight_rom[12226] = 0;
        weight_rom[12227] = -4;
        weight_rom[12228] = -2;
        weight_rom[12229] = 3;
        weight_rom[12230] = 0;
        weight_rom[12231] = -8;
        weight_rom[12232] = 10;
        weight_rom[12233] = 51;
        weight_rom[12234] = 52;
        weight_rom[12235] = 15;
        weight_rom[12236] = -1;
        weight_rom[12237] = 6;
        weight_rom[12238] = 27;
        weight_rom[12239] = 11;
        weight_rom[12240] = -3;
        weight_rom[12241] = -9;
        weight_rom[12242] = -13;
        weight_rom[12243] = 2;
        weight_rom[12244] = 7;
        weight_rom[12245] = 7;
        weight_rom[12246] = 8;
        weight_rom[12247] = 6;
        weight_rom[12248] = 32;
        weight_rom[12249] = 47;
        weight_rom[12250] = 43;
        weight_rom[12251] = 19;
        weight_rom[12252] = 8;
        weight_rom[12253] = -5;
        weight_rom[12254] = -9;
        weight_rom[12255] = 2;
        weight_rom[12256] = -10;
        weight_rom[12257] = 1;
        weight_rom[12258] = 5;
        weight_rom[12259] = 0;
        weight_rom[12260] = 3;
        weight_rom[12261] = 44;
        weight_rom[12262] = 53;
        weight_rom[12263] = 4;
        weight_rom[12264] = -4;
        weight_rom[12265] = 3;
        weight_rom[12266] = 2;
        weight_rom[12267] = 4;
        weight_rom[12268] = -9;
        weight_rom[12269] = -9;
        weight_rom[12270] = -15;
        weight_rom[12271] = -4;
        weight_rom[12272] = -4;
        weight_rom[12273] = 0;
        weight_rom[12274] = -3;
        weight_rom[12275] = 9;
        weight_rom[12276] = 34;
        weight_rom[12277] = 37;
        weight_rom[12278] = 26;
        weight_rom[12279] = 5;
        weight_rom[12280] = 8;
        weight_rom[12281] = 9;
        weight_rom[12282] = 3;
        weight_rom[12283] = 3;
        weight_rom[12284] = 6;
        weight_rom[12285] = 1;
        weight_rom[12286] = 2;
        weight_rom[12287] = 18;
        weight_rom[12288] = 21;
        weight_rom[12289] = 39;
        weight_rom[12290] = 24;
        weight_rom[12291] = 15;
        weight_rom[12292] = 1;
        weight_rom[12293] = 7;
        weight_rom[12294] = -9;
        weight_rom[12295] = 3;
        weight_rom[12296] = -6;
        weight_rom[12297] = -19;
        weight_rom[12298] = -15;
        weight_rom[12299] = -6;
        weight_rom[12300] = -13;
        weight_rom[12301] = 2;
        weight_rom[12302] = 3;
        weight_rom[12303] = 9;
        weight_rom[12304] = 4;
        weight_rom[12305] = 19;
        weight_rom[12306] = 16;
        weight_rom[12307] = 15;
        weight_rom[12308] = 15;
        weight_rom[12309] = 22;
        weight_rom[12310] = 7;
        weight_rom[12311] = -2;
        weight_rom[12312] = -5;
        weight_rom[12313] = 8;
        weight_rom[12314] = 17;
        weight_rom[12315] = 9;
        weight_rom[12316] = -9;
        weight_rom[12317] = 6;
        weight_rom[12318] = 34;
        weight_rom[12319] = 6;
        weight_rom[12320] = 3;
        weight_rom[12321] = -8;
        weight_rom[12322] = 1;
        weight_rom[12323] = 17;
        weight_rom[12324] = 17;
        weight_rom[12325] = -8;
        weight_rom[12326] = 2;
        weight_rom[12327] = 22;
        weight_rom[12328] = 0;
        weight_rom[12329] = 12;
        weight_rom[12330] = 16;
        weight_rom[12331] = 11;
        weight_rom[12332] = 20;
        weight_rom[12333] = 8;
        weight_rom[12334] = 18;
        weight_rom[12335] = 23;
        weight_rom[12336] = 12;
        weight_rom[12337] = 17;
        weight_rom[12338] = 9;
        weight_rom[12339] = 10;
        weight_rom[12340] = 18;
        weight_rom[12341] = 16;
        weight_rom[12342] = -5;
        weight_rom[12343] = 3;
        weight_rom[12344] = 12;
        weight_rom[12345] = 0;
        weight_rom[12346] = 15;
        weight_rom[12347] = 0;
        weight_rom[12348] = -3;
        weight_rom[12349] = 16;
        weight_rom[12350] = 19;
        weight_rom[12351] = 30;
        weight_rom[12352] = 7;
        weight_rom[12353] = 1;
        weight_rom[12354] = 4;
        weight_rom[12355] = 14;
        weight_rom[12356] = 13;
        weight_rom[12357] = 10;
        weight_rom[12358] = 12;
        weight_rom[12359] = 22;
        weight_rom[12360] = 13;
        weight_rom[12361] = 20;
        weight_rom[12362] = 19;
        weight_rom[12363] = 11;
        weight_rom[12364] = 3;
        weight_rom[12365] = 24;
        weight_rom[12366] = 17;
        weight_rom[12367] = 26;
        weight_rom[12368] = 8;
        weight_rom[12369] = 4;
        weight_rom[12370] = 5;
        weight_rom[12371] = 14;
        weight_rom[12372] = 5;
        weight_rom[12373] = -5;
        weight_rom[12374] = -4;
        weight_rom[12375] = -1;
        weight_rom[12376] = -3;
        weight_rom[12377] = -2;
        weight_rom[12378] = 2;
        weight_rom[12379] = 15;
        weight_rom[12380] = 13;
        weight_rom[12381] = 31;
        weight_rom[12382] = 28;
        weight_rom[12383] = 22;
        weight_rom[12384] = 17;
        weight_rom[12385] = 15;
        weight_rom[12386] = 16;
        weight_rom[12387] = 13;
        weight_rom[12388] = 9;
        weight_rom[12389] = 4;
        weight_rom[12390] = 3;
        weight_rom[12391] = 8;
        weight_rom[12392] = -3;
        weight_rom[12393] = 12;
        weight_rom[12394] = 15;
        weight_rom[12395] = 20;
        weight_rom[12396] = 21;
        weight_rom[12397] = 13;
        weight_rom[12398] = -4;
        weight_rom[12399] = -14;
        weight_rom[12400] = -3;
        weight_rom[12401] = 1;
        weight_rom[12402] = 4;
        weight_rom[12403] = -3;
        weight_rom[12404] = -1;
        weight_rom[12405] = -1;
        weight_rom[12406] = 19;
        weight_rom[12407] = -13;
        weight_rom[12408] = 15;
        weight_rom[12409] = 6;
        weight_rom[12410] = 21;
        weight_rom[12411] = 19;
        weight_rom[12412] = 21;
        weight_rom[12413] = 31;
        weight_rom[12414] = 9;
        weight_rom[12415] = 17;
        weight_rom[12416] = 11;
        weight_rom[12417] = 10;
        weight_rom[12418] = 0;
        weight_rom[12419] = 11;
        weight_rom[12420] = 13;
        weight_rom[12421] = 4;
        weight_rom[12422] = 21;
        weight_rom[12423] = 32;
        weight_rom[12424] = 26;
        weight_rom[12425] = 10;
        weight_rom[12426] = -2;
        weight_rom[12427] = -4;
        weight_rom[12428] = -22;
        weight_rom[12429] = 0;
        weight_rom[12430] = 11;
        weight_rom[12431] = -2;
        weight_rom[12432] = 3;
        weight_rom[12433] = -2;
        weight_rom[12434] = 6;
        weight_rom[12435] = -35;
        weight_rom[12436] = -8;
        weight_rom[12437] = -15;
        weight_rom[12438] = -3;
        weight_rom[12439] = -3;
        weight_rom[12440] = 1;
        weight_rom[12441] = 9;
        weight_rom[12442] = 7;
        weight_rom[12443] = 8;
        weight_rom[12444] = 8;
        weight_rom[12445] = 0;
        weight_rom[12446] = 4;
        weight_rom[12447] = -8;
        weight_rom[12448] = 7;
        weight_rom[12449] = -9;
        weight_rom[12450] = -4;
        weight_rom[12451] = -6;
        weight_rom[12452] = -15;
        weight_rom[12453] = -4;
        weight_rom[12454] = -25;
        weight_rom[12455] = -23;
        weight_rom[12456] = -3;
        weight_rom[12457] = 22;
        weight_rom[12458] = -1;
        weight_rom[12459] = 5;
        weight_rom[12460] = 0;
        weight_rom[12461] = -2;
        weight_rom[12462] = 4;
        weight_rom[12463] = -7;
        weight_rom[12464] = -26;
        weight_rom[12465] = -50;
        weight_rom[12466] = -18;
        weight_rom[12467] = -35;
        weight_rom[12468] = -36;
        weight_rom[12469] = -32;
        weight_rom[12470] = -14;
        weight_rom[12471] = -30;
        weight_rom[12472] = -36;
        weight_rom[12473] = -31;
        weight_rom[12474] = -20;
        weight_rom[12475] = -21;
        weight_rom[12476] = -28;
        weight_rom[12477] = -44;
        weight_rom[12478] = -58;
        weight_rom[12479] = -65;
        weight_rom[12480] = -51;
        weight_rom[12481] = -78;
        weight_rom[12482] = -47;
        weight_rom[12483] = -39;
        weight_rom[12484] = -16;
        weight_rom[12485] = -1;
        weight_rom[12486] = 4;
        weight_rom[12487] = -4;
        weight_rom[12488] = 0;
        weight_rom[12489] = 0;
        weight_rom[12490] = 4;
        weight_rom[12491] = 1;
        weight_rom[12492] = -28;
        weight_rom[12493] = -17;
        weight_rom[12494] = -33;
        weight_rom[12495] = -30;
        weight_rom[12496] = -56;
        weight_rom[12497] = -54;
        weight_rom[12498] = -69;
        weight_rom[12499] = -79;
        weight_rom[12500] = -77;
        weight_rom[12501] = -92;
        weight_rom[12502] = -100;
        weight_rom[12503] = -77;
        weight_rom[12504] = -88;
        weight_rom[12505] = -72;
        weight_rom[12506] = -74;
        weight_rom[12507] = -65;
        weight_rom[12508] = -74;
        weight_rom[12509] = -54;
        weight_rom[12510] = -34;
        weight_rom[12511] = -11;
        weight_rom[12512] = -1;
        weight_rom[12513] = -1;
        weight_rom[12514] = 0;
        weight_rom[12515] = 3;
        weight_rom[12516] = 0;
        weight_rom[12517] = 1;
        weight_rom[12518] = -4;
        weight_rom[12519] = 4;
        weight_rom[12520] = 1;
        weight_rom[12521] = 19;
        weight_rom[12522] = 27;
        weight_rom[12523] = -9;
        weight_rom[12524] = -17;
        weight_rom[12525] = -19;
        weight_rom[12526] = -28;
        weight_rom[12527] = -27;
        weight_rom[12528] = -26;
        weight_rom[12529] = 3;
        weight_rom[12530] = -35;
        weight_rom[12531] = -17;
        weight_rom[12532] = -14;
        weight_rom[12533] = -6;
        weight_rom[12534] = -15;
        weight_rom[12535] = -22;
        weight_rom[12536] = -9;
        weight_rom[12537] = -3;
        weight_rom[12538] = -17;
        weight_rom[12539] = 0;
        weight_rom[12540] = -1;
        weight_rom[12541] = 2;
        weight_rom[12542] = -2;
        weight_rom[12543] = -2;
        weight_rom[12544] = 127;
        weight_rom[12545] = 7;
        weight_rom[12546] = -108;
        weight_rom[12547] = 85;
        weight_rom[12548] = -81;
        weight_rom[12549] = 108;
        weight_rom[12550] = -14;
        weight_rom[12551] = -25;
        weight_rom[12552] = 77;
        weight_rom[12553] = 107;
        weight_rom[12554] = 76;
        weight_rom[12555] = 9;
        weight_rom[12556] = 107;
        weight_rom[12557] = -53;
        weight_rom[12558] = -9;
        weight_rom[12559] = -14;
        weight_rom[12560] = -81;
        weight_rom[12561] = 28;
        weight_rom[12562] = -44;
        weight_rom[12563] = -5;
        weight_rom[12564] = -3;
        weight_rom[12565] = -25;
        weight_rom[12566] = 33;
        weight_rom[12567] = -89;
        weight_rom[12568] = 22;
        weight_rom[12569] = -26;
        weight_rom[12570] = -60;
        weight_rom[12571] = 21;
        weight_rom[12572] = 34;
        weight_rom[12573] = 7;
        weight_rom[12574] = -19;
        weight_rom[12575] = -55;
        weight_rom[12576] = 26;
        weight_rom[12577] = -29;
        weight_rom[12578] = -68;
        weight_rom[12579] = 39;
        weight_rom[12580] = 29;
        weight_rom[12581] = -32;
        weight_rom[12582] = -8;
        weight_rom[12583] = 32;
        weight_rom[12584] = 41;
        weight_rom[12585] = -67;
        weight_rom[12586] = 44;
        weight_rom[12587] = -31;
        weight_rom[12588] = -14;
        weight_rom[12589] = -51;
        weight_rom[12590] = 35;
        weight_rom[12591] = 24;
        weight_rom[12592] = -29;
        weight_rom[12593] = -25;
        weight_rom[12594] = -47;
        weight_rom[12595] = -88;
        weight_rom[12596] = -40;
        weight_rom[12597] = -26;
        weight_rom[12598] = 36;
        weight_rom[12599] = -31;
        weight_rom[12600] = -42;
        weight_rom[12601] = 25;
        weight_rom[12602] = 46;
        weight_rom[12603] = 23;
        weight_rom[12604] = -19;
        weight_rom[12605] = 9;
        weight_rom[12606] = 22;
        weight_rom[12607] = 35;
        weight_rom[12608] = 0;
        weight_rom[12609] = -68;
        weight_rom[12610] = 31;
        weight_rom[12611] = -21;
        weight_rom[12612] = -28;
        weight_rom[12613] = -16;
        weight_rom[12614] = 27;
        weight_rom[12615] = 55;
        weight_rom[12616] = 27;
        weight_rom[12617] = -35;
        weight_rom[12618] = -41;
        weight_rom[12619] = 10;
        weight_rom[12620] = -32;
        weight_rom[12621] = 26;
        weight_rom[12622] = 30;
        weight_rom[12623] = 2;
        weight_rom[12624] = -45;
        weight_rom[12625] = -21;
        weight_rom[12626] = 12;
        weight_rom[12627] = 2;
        weight_rom[12628] = 21;
        weight_rom[12629] = -6;
        weight_rom[12630] = -83;
        weight_rom[12631] = 20;
        weight_rom[12632] = 11;
        weight_rom[12633] = 17;
        weight_rom[12634] = -10;
        weight_rom[12635] = -90;
        weight_rom[12636] = 64;
        weight_rom[12637] = 0;
        weight_rom[12638] = 28;
        weight_rom[12639] = 13;
        weight_rom[12640] = 42;
        weight_rom[12641] = -1;
        weight_rom[12642] = -17;
        weight_rom[12643] = 15;
        weight_rom[12644] = -75;
        weight_rom[12645] = 33;
        weight_rom[12646] = -36;
        weight_rom[12647] = 62;
        weight_rom[12648] = 0;
        weight_rom[12649] = -39;
        weight_rom[12650] = 27;
        weight_rom[12651] = 46;
        weight_rom[12652] = 12;
        weight_rom[12653] = 18;
        weight_rom[12654] = -127;
        weight_rom[12655] = -52;
        weight_rom[12656] = -62;
        weight_rom[12657] = 47;
        weight_rom[12658] = -55;
        weight_rom[12659] = 47;
        weight_rom[12660] = -46;
        weight_rom[12661] = -70;
        weight_rom[12662] = -64;
        weight_rom[12663] = -30;
        weight_rom[12664] = 20;
        weight_rom[12665] = 16;
        weight_rom[12666] = 7;
        weight_rom[12667] = 11;
        weight_rom[12668] = -46;
        weight_rom[12669] = 9;
        weight_rom[12670] = -34;
        weight_rom[12671] = 26;
        weight_rom[12672] = 45;
        weight_rom[12673] = -29;
        weight_rom[12674] = 8;
        weight_rom[12675] = -23;
        weight_rom[12676] = 1;
        weight_rom[12677] = 50;
        weight_rom[12678] = 30;
        weight_rom[12679] = -79;
        weight_rom[12680] = 70;
        weight_rom[12681] = 21;
        weight_rom[12682] = -66;
        weight_rom[12683] = -37;
        weight_rom[12684] = -8;
        weight_rom[12685] = -72;
        weight_rom[12686] = 24;
        weight_rom[12687] = -3;
        weight_rom[12688] = -2;
        weight_rom[12689] = 25;
        weight_rom[12690] = 20;
        weight_rom[12691] = -33;
        weight_rom[12692] = 34;
        weight_rom[12693] = 22;
        weight_rom[12694] = -19;
        weight_rom[12695] = -24;
        weight_rom[12696] = -66;
        weight_rom[12697] = -67;
        weight_rom[12698] = 11;
        weight_rom[12699] = 17;
        weight_rom[12700] = -30;
        weight_rom[12701] = 24;
        weight_rom[12702] = -38;
        weight_rom[12703] = 2;
        weight_rom[12704] = -14;
        weight_rom[12705] = 21;
        weight_rom[12706] = 36;
        weight_rom[12707] = -32;
        weight_rom[12708] = 53;
        weight_rom[12709] = -20;
        weight_rom[12710] = 17;
        weight_rom[12711] = 56;
        weight_rom[12712] = -38;
        weight_rom[12713] = 21;
        weight_rom[12714] = 18;
        weight_rom[12715] = -52;
        weight_rom[12716] = 9;
        weight_rom[12717] = -45;
        weight_rom[12718] = -11;
        weight_rom[12719] = -48;
        weight_rom[12720] = -2;
        weight_rom[12721] = 88;
        weight_rom[12722] = 16;
        weight_rom[12723] = -44;
        weight_rom[12724] = 11;
        weight_rom[12725] = 95;
        weight_rom[12726] = -34;
        weight_rom[12727] = 0;
        weight_rom[12728] = -127;
        weight_rom[12729] = -46;
    end

    // 主状态机和MAC单元
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            valid <= 0;
            digit_out <= 0;
            neuron_idx <= 0;
            input_idx <= 0;
            accumulator <= 0;
        end else begin
            case (state)
                IDLE: begin
                    valid <= 0;
                    digit_out <= 0;
                    neuron_idx <= 0;
                    input_idx <= 0;
                    if (start) begin
                        state <= LAYER1_COMPUTE;
                        // 初始化累加器为第一个神经元的偏置 (地址12544)
                        accumulator <= $signed(weight_rom[12544]);
                    end
                end

                LAYER1_COMPUTE: begin
                    // MAC操作: accumulator += weight * input
                    // 读取Layer1权重: 地址 = neuron_idx * 784 + input_idx
                    accumulator <= accumulator + ($signed(weight_rom[neuron_idx * 784 + input_idx]) * $signed({31'b0, image_in[input_idx]}));

                    if (input_idx == 783) begin
                        // 当前神经元计算完成，进入激活
                        state <= LAYER1_ACTIVATE;
                        input_idx <= 0;
                    end else begin
                        // 继续计算下一个输入
                        input_idx <= input_idx + 1;
                    end
                end

                LAYER1_ACTIVATE: begin
                    // ReLU激活
                    if (accumulator < 0) begin
                        layer1_out[neuron_idx] <= 0;
                    end else begin
                        layer1_out[neuron_idx] <= accumulator;
                    end

                    if (neuron_idx == 15) begin
                        // Layer1完成，进入Layer2
                        state <= LAYER2_COMPUTE;
                        neuron_idx <= 0;
                        input_idx <= 0;
                        // 初始化为Layer2第一个神经元的偏置 (地址12720)
                        accumulator <= $signed(weight_rom[12720]);
                    end else begin
                        // 计算下一个神经元
                        neuron_idx <= neuron_idx + 1;
                        input_idx <= 0;
                        state <= LAYER1_COMPUTE;
                        // 加载下一个神经元的偏置 (地址 12544 + neuron_idx + 1)
                        accumulator <= $signed(weight_rom[12544 + neuron_idx + 1]);
                    end
                end

                LAYER2_COMPUTE: begin
                    // MAC操作: accumulator += (weight * layer1_out) >> 7
                    // 读取Layer2权重: 地址 = 12560 + neuron_idx * 16 + input_idx
                    accumulator <= accumulator + (($signed(weight_rom[12560 + neuron_idx * 16 + input_idx]) * layer1_out[input_idx]) >>> 7);

                    if (input_idx == 15) begin
                        // 当前神经元计算完成
                        layer2_out[neuron_idx] <= accumulator;

                        if (neuron_idx == 9) begin
                            // Layer2完成，进入argmax
                            state <= ARGMAX;
                        end else begin
                            // 计算下一个神经元
                            neuron_idx <= neuron_idx + 1;
                            input_idx <= 0;
                            // 加载下一个神经元的偏置 (地址 12720 + neuron_idx + 1)
                            accumulator <= $signed(weight_rom[12720 + neuron_idx + 1]);
                        end
                    end else begin
                        // 继续计算下一个输入
                        input_idx <= input_idx + 1;
                    end
                end

                ARGMAX: begin
                    // 找到最大值的索引（使用串行比较减少组合逻辑）
                    if (layer2_out[0] >= layer2_out[1] && layer2_out[0] >= layer2_out[2] &&
                        layer2_out[0] >= layer2_out[3] && layer2_out[0] >= layer2_out[4] &&
                        layer2_out[0] >= layer2_out[5] && layer2_out[0] >= layer2_out[6] &&
                        layer2_out[0] >= layer2_out[7] && layer2_out[0] >= layer2_out[8] &&
                        layer2_out[0] >= layer2_out[9])
                        digit_out <= 0;
                    else if (layer2_out[1] >= layer2_out[2] && layer2_out[1] >= layer2_out[3] &&
                             layer2_out[1] >= layer2_out[4] && layer2_out[1] >= layer2_out[5] &&
                             layer2_out[1] >= layer2_out[6] && layer2_out[1] >= layer2_out[7] &&
                             layer2_out[1] >= layer2_out[8] && layer2_out[1] >= layer2_out[9])
                        digit_out <= 1;
                    else if (layer2_out[2] >= layer2_out[3] && layer2_out[2] >= layer2_out[4] &&
                             layer2_out[2] >= layer2_out[5] && layer2_out[2] >= layer2_out[6] &&
                             layer2_out[2] >= layer2_out[7] && layer2_out[2] >= layer2_out[8] &&
                             layer2_out[2] >= layer2_out[9])
                        digit_out <= 2;
                    else if (layer2_out[3] >= layer2_out[4] && layer2_out[3] >= layer2_out[5] &&
                             layer2_out[3] >= layer2_out[6] && layer2_out[3] >= layer2_out[7] &&
                             layer2_out[3] >= layer2_out[8] && layer2_out[3] >= layer2_out[9])
                        digit_out <= 3;
                    else if (layer2_out[4] >= layer2_out[5] && layer2_out[4] >= layer2_out[6] &&
                             layer2_out[4] >= layer2_out[7] && layer2_out[4] >= layer2_out[8] &&
                             layer2_out[4] >= layer2_out[9])
                        digit_out <= 4;
                    else if (layer2_out[5] >= layer2_out[6] && layer2_out[5] >= layer2_out[7] &&
                             layer2_out[5] >= layer2_out[8] && layer2_out[5] >= layer2_out[9])
                        digit_out <= 5;
                    else if (layer2_out[6] >= layer2_out[7] && layer2_out[6] >= layer2_out[8] &&
                             layer2_out[6] >= layer2_out[9])
                        digit_out <= 6;
                    else if (layer2_out[7] >= layer2_out[8] && layer2_out[7] >= layer2_out[9])
                        digit_out <= 7;
                    else if (layer2_out[8] >= layer2_out[9])
                        digit_out <= 8;
                    else
                        digit_out <= 9;

                    valid <= 1;
                    state <= DONE;
                end

                DONE: begin
                    // 保持结果直到下一次start
                    valid <= 1;
                    // 允许在DONE状态重新开始新的计算
                    if (start) begin
                        state <= LAYER1_COMPUTE;
                        neuron_idx <= 0;
                        input_idx <= 0;
                        valid <= 0;
                        digit_out <= 0;
                        // 初始化累加器为第一个神经元的偏置 (地址12544)
                        accumulator <= $signed(weight_rom[12544]);
                    end
                end

                default: begin
                    state <= IDLE;
                end
            endcase
        end
    end

endmodule
