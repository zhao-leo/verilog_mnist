// MNIST手写数字识别模型 - Int8量化版本
// 输入: 28x28二值图像 (784位)
// 输出: 预测数字 (0-9)

module mnist_model(
    input wire clk,
    input wire rst,
    input wire [783:0] image_in,  // 28*28 = 784位输入
    input wire start,
    output reg [3:0] digit_out,   // 输出数字 0-9
    output reg valid
);

    // 状态机
    localparam IDLE = 2'd0;
    localparam LAYER1 = 2'd1;
    localparam LAYER2 = 2'd2;
    localparam DONE = 2'd3;

    reg [1:0] state;
    reg [9:0] counter;

    // 第一层输出 (16个神经元)
    reg signed [31:0] layer1_out [0:15];

    // 第二层输出 (10个神经元)
    reg signed [31:0] layer2_out [0:9];

    integer i;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            valid <= 0;
            digit_out <= 0;
            counter <= 0;
        end else begin
            case (state)
                IDLE: begin
                    valid <= 0;
                    if (start) begin
                        state <= LAYER1;
                        counter <= 0;
                    end
                end

                LAYER1: begin
                    // 计算第一层（简化：直接计算所有神经元）
                    if (counter == 0) begin
                        layer1_out[0] = 75 -3 * image_in[0] -1 * image_in[1] +5 * image_in[2] +4 * image_in[3] +1 * image_in[4] -1 * image_in[5] +4 * image_in[6] -6 * image_in[7] -2 * image_in[8] -1 * image_in[9] -2 * image_in[10] -5 * image_in[11] -4 * image_in[12] -5 * image_in[13] +8 * image_in[14] +1 * image_in[15] +6 * image_in[16] -1 * image_in[17] +1 * image_in[18] +1 * image_in[19] -1 * image_in[20] -2 * image_in[22] -2 * image_in[23] +1 * image_in[24] +3 * image_in[25] -5 * image_in[26] -3 * image_in[27] +3 * image_in[28] -6 * image_in[29] +5 * image_in[30] -1 * image_in[31]
                            +1 * image_in[32] +2 * image_in[33] -13 * image_in[34] -20 * image_in[35] -11 * image_in[36] -16 * image_in[37] -27 * image_in[38] -17 * image_in[39] -39 * image_in[40] -52 * image_in[41] +14 * image_in[42] +6 * image_in[43] +25 * image_in[44] -15 * image_in[45] -42 * image_in[46] -26 * image_in[47] -22 * image_in[48] -13 * image_in[49] -24 * image_in[50] -15 * image_in[51] -5 * image_in[53] +2 * image_in[54] +2 * image_in[55] -5 * image_in[56] -1 * image_in[57] -1 * image_in[59] -14 * image_in[60] -4 * image_in[61] -12 * image_in[62] -36 * image_in[63]
                            -36 * image_in[64] -12 * image_in[65] -40 * image_in[66] -25 * image_in[67] -27 * image_in[68] -13 * image_in[69] -20 * image_in[70] +1 * image_in[71] -6 * image_in[72] -11 * image_in[73] -15 * image_in[74] -22 * image_in[75] -55 * image_in[76] -33 * image_in[77] -36 * image_in[78] -26 * image_in[79] -7 * image_in[80] +16 * image_in[81] +3 * image_in[82] -2 * image_in[83] -5 * image_in[85] -11 * image_in[86] -2 * image_in[87] -4 * image_in[88] -32 * image_in[89] -21 * image_in[90] -25 * image_in[91] -27 * image_in[92] -14 * image_in[93] -25 * image_in[94] -35 * image_in[95]
                            -23 * image_in[96] -14 * image_in[97] -13 * image_in[98] -14 * image_in[99] +2 * image_in[100] -8 * image_in[101] -25 * image_in[102] -26 * image_in[103] -15 * image_in[104] +3 * image_in[105] -15 * image_in[106] -17 * image_in[107] -27 * image_in[108] +35 * image_in[109] -1 * image_in[111] +2 * image_in[112] -5 * image_in[113] +18 * image_in[114] -5 * image_in[115] -34 * image_in[116] -35 * image_in[117] -5 * image_in[118] -12 * image_in[119] -17 * image_in[120] +3 * image_in[121] +6 * image_in[122] +27 * image_in[123] +24 * image_in[124] +14 * image_in[125] +33 * image_in[126] +30 * image_in[127]
                            +27 * image_in[128] +17 * image_in[129] +14 * image_in[130] +2 * image_in[131] +1 * image_in[132] +19 * image_in[133] -3 * image_in[134] +11 * image_in[135] +41 * image_in[136] +25 * image_in[137] +26 * image_in[138] +6 * image_in[139] +5 * image_in[140] +6 * image_in[142] -11 * image_in[143] -42 * image_in[144] -31 * image_in[145] -23 * image_in[146] -13 * image_in[147] -14 * image_in[148] +2 * image_in[149] +5 * image_in[150] +21 * image_in[151] +19 * image_in[152] +14 * image_in[153] +12 * image_in[154] +16 * image_in[155] +28 * image_in[156] +32 * image_in[157] +14 * image_in[158] +17 * image_in[159]
                            +35 * image_in[160] +29 * image_in[161] +28 * image_in[162] +22 * image_in[163] +18 * image_in[164] +39 * image_in[165] -1 * image_in[168] +5 * image_in[169] -31 * image_in[170] -48 * image_in[171] -46 * image_in[172] -8 * image_in[173] -18 * image_in[174] -12 * image_in[175] -11 * image_in[176] -6 * image_in[177] +1 * image_in[178] +8 * image_in[179] +16 * image_in[180] +9 * image_in[181] +11 * image_in[182] +15 * image_in[183] +9 * image_in[184] +13 * image_in[185] +13 * image_in[186] +28 * image_in[187] +25 * image_in[188] +19 * image_in[189] +19 * image_in[190] +27 * image_in[191]
                            +58 * image_in[192] +55 * image_in[193] +33 * image_in[194] -5 * image_in[196] -32 * image_in[197] -6 * image_in[198] -62 * image_in[199] -28 * image_in[200] -25 * image_in[201] -15 * image_in[202] -22 * image_in[203] +14 * image_in[204] -8 * image_in[205] +9 * image_in[206] +3 * image_in[207] -7 * image_in[208] +3 * image_in[209] -7 * image_in[210] -1 * image_in[211] +19 * image_in[212] +16 * image_in[214] +25 * image_in[215] +25 * image_in[216] +20 * image_in[217] +32 * image_in[218] +40 * image_in[219] +49 * image_in[220] +70 * image_in[221] +16 * image_in[222] +8 * image_in[223]
                            -13 * image_in[224] -25 * image_in[225] -11 * image_in[226] -34 * image_in[227] -46 * image_in[228] -30 * image_in[229] -5 * image_in[230] -4 * image_in[231] -8 * image_in[232] +11 * image_in[233] +16 * image_in[234] +11 * image_in[235] +13 * image_in[236] +13 * image_in[237] +1 * image_in[238] -5 * image_in[239] -7 * image_in[240] +23 * image_in[242] +19 * image_in[243] +19 * image_in[244] +16 * image_in[245] +24 * image_in[246] +60 * image_in[247] +86 * image_in[248] +102 * image_in[249] +76 * image_in[250] +35 * image_in[251] -7 * image_in[252] -27 * image_in[253] -19 * image_in[254] -56 * image_in[255]
                            -53 * image_in[256] -4 * image_in[257] -4 * image_in[258] -18 * image_in[259] +8 * image_in[260] +20 * image_in[261] +23 * image_in[262] +50 * image_in[263] +42 * image_in[264] +20 * image_in[265] -13 * image_in[266] -25 * image_in[267] -5 * image_in[268] +1 * image_in[269] +12 * image_in[270] +9 * image_in[271] +11 * image_in[272] +8 * image_in[273] +16 * image_in[274] +52 * image_in[275] +94 * image_in[276] +114 * image_in[277] +48 * image_in[278] -15 * image_in[279] -9 * image_in[280] -17 * image_in[281] -12 * image_in[282] -50 * image_in[283] -9 * image_in[284] -5 * image_in[285] -1 * image_in[286] +4 * image_in[287]
                            +21 * image_in[288] +45 * image_in[289] +38 * image_in[290] +48 * image_in[291] +47 * image_in[292] -6 * image_in[293] -16 * image_in[294] -16 * image_in[295] -24 * image_in[296] -7 * image_in[297] -13 * image_in[298] -5 * image_in[299] -20 * image_in[300] +1 * image_in[301] -5 * image_in[302] +21 * image_in[303] +76 * image_in[304] +103 * image_in[305] +62 * image_in[306] +21 * image_in[307] -11 * image_in[308] -24 * image_in[309] -39 * image_in[310] -69 * image_in[311] -11 * image_in[312] +13 * image_in[313] +21 * image_in[314] +3 * image_in[315] +30 * image_in[316] +22 * image_in[317] +19 * image_in[318] +11 * image_in[319]
                            +7 * image_in[320] -1 * image_in[321] -8 * image_in[322] -3 * image_in[323] -16 * image_in[324] -10 * image_in[325] -7 * image_in[326] -8 * image_in[327] -36 * image_in[328] -22 * image_in[329] -17 * image_in[330] +1 * image_in[331] +56 * image_in[332] +81 * image_in[333] +73 * image_in[334] -13 * image_in[335] -13 * image_in[336] -13 * image_in[337] -18 * image_in[338] -20 * image_in[339] +17 * image_in[340] +11 * image_in[341] +14 * image_in[342] +6 * image_in[343] +8 * image_in[344] +7 * image_in[345] +13 * image_in[346] +5 * image_in[347] +2 * image_in[348] +16 * image_in[349] +10 * image_in[350] -1 * image_in[351]
                            -18 * image_in[352] -23 * image_in[353] -20 * image_in[354] +7 * image_in[355] +5 * image_in[356] -7 * image_in[357] -43 * image_in[358] -49 * image_in[359] -9 * image_in[360] +47 * image_in[361] +63 * image_in[362] -17 * image_in[363] -6 * image_in[364] +1 * image_in[365] -40 * image_in[366] -4 * image_in[367] +4 * image_in[368] -4 * image_in[369] -20 * image_in[370] -10 * image_in[371] +8 * image_in[372] +6 * image_in[373] +7 * image_in[374] +20 * image_in[375] +44 * image_in[376] +28 * image_in[377] +15 * image_in[378] +15 * image_in[379] -18 * image_in[380] -17 * image_in[381] -11 * image_in[382] +4 * image_in[383]
                            +16 * image_in[384] -23 * image_in[385] -18 * image_in[386] -37 * image_in[387] -20 * image_in[388] +39 * image_in[389] +78 * image_in[390] +35 * image_in[391] -4 * image_in[392] -16 * image_in[393] -15 * image_in[394] -21 * image_in[395] +7 * image_in[396] -9 * image_in[397] -11 * image_in[398] +3 * image_in[399] +3 * image_in[400] +21 * image_in[401] +21 * image_in[402] +22 * image_in[403] +34 * image_in[404] +49 * image_in[405] +40 * image_in[406] +20 * image_in[407] -2 * image_in[408] -8 * image_in[409] -18 * image_in[410] -19 * image_in[411] -11 * image_in[412] -23 * image_in[413] -24 * image_in[414] -29 * image_in[415]
                            -1 * image_in[416] +14 * image_in[417] +50 * image_in[418] -2 * image_in[419] +1 * image_in[420] -14 * image_in[421] -41 * image_in[422] +15 * image_in[423] +5 * image_in[424] -17 * image_in[425] -7 * image_in[426] -4 * image_in[427] +27 * image_in[428] +22 * image_in[429] +17 * image_in[430] +15 * image_in[431] +33 * image_in[432] +48 * image_in[433] +37 * image_in[434] +21 * image_in[435] +16 * image_in[436] -9 * image_in[437] -10 * image_in[438] -24 * image_in[439] -51 * image_in[440] -43 * image_in[441] -35 * image_in[442] -33 * image_in[443] +28 * image_in[445] +51 * image_in[446] +11 * image_in[447]
                            +4 * image_in[448] -1 * image_in[449] -32 * image_in[450] +42 * image_in[451] -4 * image_in[452] -7 * image_in[453] +10 * image_in[454] -11 * image_in[455] -5 * image_in[456] +6 * image_in[458] +9 * image_in[459] +37 * image_in[460] +40 * image_in[461] +37 * image_in[462] +26 * image_in[463] +11 * image_in[464] -2 * image_in[465] -24 * image_in[466] -35 * image_in[467] -35 * image_in[468] -22 * image_in[469] -6 * image_in[470] -1 * image_in[471] +14 * image_in[472] +52 * image_in[473] +80 * image_in[474] +30 * image_in[475] -3 * image_in[476] -14 * image_in[477] +7 * image_in[478] +17 * image_in[479] +14 * image_in[481] +35 * image_in[482] +9 * image_in[483] +2 * image_in[484] +9 * image_in[485] +11 * image_in[486] +5 * image_in[487] +26 * image_in[488] +30 * image_in[489] +27 * image_in[490] +22 * image_in[491] +23 * image_in[492] -1 * image_in[493] -9 * image_in[494] -20 * image_in[495] -6 * image_in[496] -5 * image_in[497] -7 * image_in[498] +47 * image_in[500] +30 * image_in[501] +79 * image_in[502] -4 * image_in[503] -12 * image_in[505] -9 * image_in[506] -7 * image_in[507] +21 * image_in[508] +49 * image_in[509] +46 * image_in[510] +28 * image_in[511]
                            +25 * image_in[512] +7 * image_in[513] +5 * image_in[514] +13 * image_in[515] +22 * image_in[516] +33 * image_in[517] +28 * image_in[518] +11 * image_in[519] -1 * image_in[520] -12 * image_in[521] -15 * image_in[522] -1 * image_in[523] +17 * image_in[524] +18 * image_in[526] +38 * image_in[527] +77 * image_in[528] +28 * image_in[529] +22 * image_in[530] +30 * image_in[531] -1 * image_in[532] -12 * image_in[533] +12 * image_in[534] -21 * image_in[535] +26 * image_in[536] +35 * image_in[537] +29 * image_in[538] +32 * image_in[539] +32 * image_in[540] +14 * image_in[541] +6 * image_in[542] +2 * image_in[543]
                            -5 * image_in[544] +27 * image_in[545] +1 * image_in[546] +8 * image_in[547] -2 * image_in[548] -5 * image_in[549] +7 * image_in[550] +10 * image_in[551] +15 * image_in[552] +3 * image_in[553] +32 * image_in[554] +54 * image_in[555] +56 * image_in[556] +56 * image_in[557] +30 * image_in[558] +14 * image_in[559] -8 * image_in[561] +8 * image_in[562] -14 * image_in[563] +3 * image_in[564] +18 * image_in[565] +32 * image_in[566] +20 * image_in[567] +18 * image_in[568] +19 * image_in[569] +12 * image_in[570] -2 * image_in[571] -10 * image_in[572] -3 * image_in[573] -20 * image_in[574] -8 * image_in[575]
                            +4 * image_in[576] +16 * image_in[577] +21 * image_in[578] +13 * image_in[579] +21 * image_in[580] +45 * image_in[581] +75 * image_in[582] +66 * image_in[583] +50 * image_in[584] +26 * image_in[585] +11 * image_in[586] +3 * image_in[587] +3 * image_in[588] -15 * image_in[589] +1 * image_in[590] -7 * image_in[591] +17 * image_in[592] +26 * image_in[593] +37 * image_in[594] +26 * image_in[595] +24 * image_in[596] +26 * image_in[597] -4 * image_in[598] +6 * image_in[599] -3 * image_in[600] -7 * image_in[601] -4 * image_in[602] +4 * image_in[603] -3 * image_in[604] +8 * image_in[605] +10 * image_in[606] +25 * image_in[607]
                            +37 * image_in[608] +53 * image_in[609] +66 * image_in[610] +99 * image_in[611] +48 * image_in[612] +32 * image_in[613] -1 * image_in[614] +4 * image_in[615] -6 * image_in[617] -6 * image_in[618] -10 * image_in[619] +19 * image_in[620] +17 * image_in[621] +23 * image_in[622] +31 * image_in[623] +17 * image_in[624] +7 * image_in[625] +12 * image_in[626] +9 * image_in[627] +3 * image_in[628] +6 * image_in[629] +6 * image_in[630] +3 * image_in[631] +4 * image_in[632] +12 * image_in[633] +32 * image_in[634] +22 * image_in[635] +37 * image_in[636] +56 * image_in[637] +54 * image_in[638] +59 * image_in[639]
                            +41 * image_in[640] +19 * image_in[641] +1 * image_in[642] +2 * image_in[643] -4 * image_in[644] +5 * image_in[645] -9 * image_in[646] -18 * image_in[647] -12 * image_in[648] -9 * image_in[649] -14 * image_in[650] -12 * image_in[651] +28 * image_in[652] +31 * image_in[653] +25 * image_in[654] +29 * image_in[655] +35 * image_in[656] +29 * image_in[657] +12 * image_in[658] +7 * image_in[659] +30 * image_in[660] +20 * image_in[661] +11 * image_in[662] +39 * image_in[663] +51 * image_in[664] +42 * image_in[665] +48 * image_in[666] +59 * image_in[667] +24 * image_in[668] +37 * image_in[669] -22 * image_in[670] +2 * image_in[671]
                            -1 * image_in[672] -2 * image_in[673] +7 * image_in[674] -40 * image_in[675] -56 * image_in[676] -62 * image_in[677] -41 * image_in[678] -41 * image_in[679] -9 * image_in[680] +24 * image_in[681] -2 * image_in[682] +16 * image_in[683] +30 * image_in[684] +23 * image_in[685] +23 * image_in[686] +25 * image_in[687] +7 * image_in[688] +11 * image_in[689] +40 * image_in[690] +31 * image_in[691] +22 * image_in[692] +23 * image_in[693] +11 * image_in[694] +26 * image_in[695] +32 * image_in[696] +39 * image_in[697] -2 * image_in[698] -3 * image_in[699] +1 * image_in[701] +9 * image_in[703]
                            -28 * image_in[704] -61 * image_in[705] -29 * image_in[706] -55 * image_in[707] -58 * image_in[708] -51 * image_in[709] -29 * image_in[710] -37 * image_in[711] -22 * image_in[712] -19 * image_in[713] -16 * image_in[714] -8 * image_in[715] +3 * image_in[716] +11 * image_in[717] -12 * image_in[718] -23 * image_in[719] -17 * image_in[720] -25 * image_in[721] +8 * image_in[722] +16 * image_in[723] +10 * image_in[724] +2 * image_in[725] +2 * image_in[726] -2 * image_in[727] +1 * image_in[728] -2 * image_in[729] -2 * image_in[730] +3 * image_in[731] -26 * image_in[732] -15 * image_in[733] -22 * image_in[734] -60 * image_in[735]
                            -77 * image_in[736] -52 * image_in[737] -49 * image_in[738] -42 * image_in[739] -24 * image_in[740] -48 * image_in[741] -61 * image_in[742] -33 * image_in[743] -47 * image_in[744] -56 * image_in[745] -56 * image_in[746] -67 * image_in[747] -21 * image_in[748] -24 * image_in[749] -16 * image_in[750] -20 * image_in[751] +2 * image_in[752] -1 * image_in[753] +4 * image_in[755] +3 * image_in[756] +1 * image_in[757] +4 * image_in[758] +1 * image_in[759] -5 * image_in[760] -17 * image_in[761] -28 * image_in[762] -34 * image_in[763] -36 * image_in[764] -23 * image_in[765] -44 * image_in[766] -7 * image_in[767]
                            -14 * image_in[768] -40 * image_in[769] -37 * image_in[770] -15 * image_in[771] -10 * image_in[772] -44 * image_in[773] -63 * image_in[774] -10 * image_in[775] -9 * image_in[776] -16 * image_in[777] -9 * image_in[778] -1 * image_in[779] -2 * image_in[780] -2 * image_in[781] +5 * image_in[782] +6 * image_in[783];
                        if (layer1_out[0] < 0) layer1_out[0] = 0;
                        layer1_out[1] = -74 -4 * image_in[0] -4 * image_in[1] -3 * image_in[2] +4 * image_in[3] -5 * image_in[4] -2 * image_in[5] +3 * image_in[6] -2 * image_in[7] +1 * image_in[8] -2 * image_in[9] +3 * image_in[10] -1 * image_in[11] -1 * image_in[12] +12 * image_in[13] +11 * image_in[14] -1 * image_in[15] +3 * image_in[16] -1 * image_in[17] +4 * image_in[18] +3 * image_in[19] -4 * image_in[20] -2 * image_in[21] -2 * image_in[22] -2 * image_in[23] +4 * image_in[24] +5 * image_in[25] -6 * image_in[26] -1 * image_in[27] +3 * image_in[28] +2 * image_in[29] +4 * image_in[30] -4 * image_in[31]
                            -5 * image_in[32] +3 * image_in[33] +12 * image_in[34] +15 * image_in[35] +11 * image_in[36] -5 * image_in[37] -1 * image_in[38] -3 * image_in[39] -18 * image_in[41] +6 * image_in[42] +18 * image_in[43] +51 * image_in[44] +8 * image_in[45] -26 * image_in[46] -23 * image_in[47] -18 * image_in[48] +7 * image_in[49] +5 * image_in[50] +1 * image_in[51] -6 * image_in[52] -6 * image_in[53] +3 * image_in[54] -5 * image_in[55] -5 * image_in[56] -5 * image_in[57] +6 * image_in[59] -13 * image_in[60] +1 * image_in[61] -5 * image_in[62] -9 * image_in[63]
                            +2 * image_in[64] +17 * image_in[65] -18 * image_in[66] +10 * image_in[67] +15 * image_in[68] +38 * image_in[69] +27 * image_in[70] +3 * image_in[71] +27 * image_in[72] -2 * image_in[73] -26 * image_in[74] -37 * image_in[75] -37 * image_in[76] -22 * image_in[77] -47 * image_in[78] -7 * image_in[79] +11 * image_in[80] +11 * image_in[81] -5 * image_in[82] -1 * image_in[83] +4 * image_in[84] +2 * image_in[86] +4 * image_in[87] -3 * image_in[88] +35 * image_in[89] +8 * image_in[90] +23 * image_in[91] +53 * image_in[92] +34 * image_in[93] +46 * image_in[94] +69 * image_in[95]
                            +83 * image_in[96] +73 * image_in[97] +78 * image_in[98] +46 * image_in[99] +34 * image_in[100] +32 * image_in[101] +21 * image_in[102] -8 * image_in[103] -7 * image_in[104] -47 * image_in[105] -60 * image_in[106] -42 * image_in[107] -13 * image_in[108] +8 * image_in[109] -4 * image_in[110] +2 * image_in[111] -3 * image_in[112] +1 * image_in[113] +18 * image_in[114] +5 * image_in[115] -2 * image_in[116] +39 * image_in[117] +25 * image_in[118] +28 * image_in[119] +44 * image_in[120] +47 * image_in[121] +58 * image_in[122] +46 * image_in[123] +51 * image_in[124] +51 * image_in[125] +52 * image_in[126] +45 * image_in[127]
                            +28 * image_in[128] +19 * image_in[129] +33 * image_in[130] +12 * image_in[131] -3 * image_in[132] -40 * image_in[133] -37 * image_in[134] -70 * image_in[135] -68 * image_in[136] -17 * image_in[137] +2 * image_in[138] +2 * image_in[139] -6 * image_in[140] +5 * image_in[141] -5 * image_in[142] +21 * image_in[143] +31 * image_in[144] +20 * image_in[145] +21 * image_in[146] +27 * image_in[147] +9 * image_in[148] +17 * image_in[149] +20 * image_in[150] +14 * image_in[151] +28 * image_in[152] +29 * image_in[153] +29 * image_in[154] +41 * image_in[155] +34 * image_in[156] +22 * image_in[157] +17 * image_in[158] +12 * image_in[159]
                            +4 * image_in[160] -16 * image_in[161] -11 * image_in[162] -44 * image_in[163] -55 * image_in[164] -9 * image_in[165] -14 * image_in[166] -2 * image_in[167] +5 * image_in[168] -1 * image_in[169] +18 * image_in[170] +46 * image_in[171] +39 * image_in[172] +8 * image_in[173] +26 * image_in[174] +1 * image_in[175] +17 * image_in[176] +13 * image_in[177] +14 * image_in[178] +14 * image_in[179] +16 * image_in[180] +36 * image_in[181] +29 * image_in[182] +36 * image_in[183] +31 * image_in[184] +19 * image_in[185] +25 * image_in[186] +6 * image_in[187] +5 * image_in[188] -5 * image_in[189] -8 * image_in[190] -25 * image_in[191]
                            -49 * image_in[192] -20 * image_in[193] -29 * image_in[194] -31 * image_in[195] +1 * image_in[196] +29 * image_in[197] +10 * image_in[198] +58 * image_in[199] +50 * image_in[200] +27 * image_in[201] +21 * image_in[202] +11 * image_in[203] +17 * image_in[204] +8 * image_in[205] +13 * image_in[206] +13 * image_in[207] +28 * image_in[208] +33 * image_in[209] +37 * image_in[210] +34 * image_in[211] +21 * image_in[212] +28 * image_in[213] +16 * image_in[214] +28 * image_in[215] +2 * image_in[216] +9 * image_in[217] +4 * image_in[218] -26 * image_in[219] -57 * image_in[220] -42 * image_in[221] -18 * image_in[222] +3 * image_in[223]
                            -1 * image_in[224] +10 * image_in[225] +17 * image_in[226] +41 * image_in[227] +62 * image_in[228] +18 * image_in[229] +16 * image_in[230] +18 * image_in[231] +4 * image_in[232] +7 * image_in[233] +22 * image_in[234] +14 * image_in[235] +33 * image_in[236] +32 * image_in[237] +42 * image_in[238] +33 * image_in[239] +44 * image_in[240] +46 * image_in[241] +37 * image_in[242] +33 * image_in[243] +32 * image_in[244] +12 * image_in[245] +34 * image_in[246] -27 * image_in[247] -87 * image_in[248] -56 * image_in[249] -9 * image_in[250] -13 * image_in[251] +1 * image_in[252] +13 * image_in[253] +8 * image_in[254] +46 * image_in[255]
                            +61 * image_in[256] +31 * image_in[257] -6 * image_in[258] -1 * image_in[259] -12 * image_in[260] +3 * image_in[261] -19 * image_in[262] -26 * image_in[263] -32 * image_in[264] -17 * image_in[265] +12 * image_in[266] +26 * image_in[267] +27 * image_in[268] +47 * image_in[269] +38 * image_in[270] +42 * image_in[271] +38 * image_in[272] +19 * image_in[273] +34 * image_in[274] -31 * image_in[275] -83 * image_in[276] -41 * image_in[277] -5 * image_in[278] +7 * image_in[279] +12 * image_in[280] +1 * image_in[281] +10 * image_in[282] +41 * image_in[283] +11 * image_in[284] -7 * image_in[285] -7 * image_in[286] -39 * image_in[287]
                            -54 * image_in[288] -61 * image_in[289] -63 * image_in[290] -68 * image_in[291] -79 * image_in[292] -56 * image_in[293] -15 * image_in[294] -6 * image_in[295] +20 * image_in[296] +29 * image_in[297] +29 * image_in[298] +28 * image_in[299] +39 * image_in[300] +38 * image_in[301] +20 * image_in[302] -27 * image_in[303] -52 * image_in[304] -42 * image_in[305] -31 * image_in[306] -8 * image_in[307] +6 * image_in[308] +10 * image_in[309] +8 * image_in[310] +20 * image_in[311] -18 * image_in[312] -56 * image_in[313] -73 * image_in[314] -72 * image_in[315] -68 * image_in[316] -62 * image_in[317] -66 * image_in[318] -57 * image_in[319]
                            -72 * image_in[320] -54 * image_in[321] -20 * image_in[322] -21 * image_in[323] -22 * image_in[324] +2 * image_in[325] +13 * image_in[326] +34 * image_in[327] +36 * image_in[328] +16 * image_in[329] +35 * image_in[330] +4 * image_in[331] -23 * image_in[332] +3 * image_in[333] +4 * image_in[334] -6 * image_in[335] +5 * image_in[336] +3 * image_in[337] -9 * image_in[338] -11 * image_in[339] -64 * image_in[340] -90 * image_in[341] -101 * image_in[342] -75 * image_in[343] -57 * image_in[344] -34 * image_in[345] -26 * image_in[346] -45 * image_in[347] -37 * image_in[348] -34 * image_in[349] -16 * image_in[350] -13 * image_in[351]
                            -4 * image_in[352] -9 * image_in[353] +5 * image_in[354] +10 * image_in[355] +18 * image_in[356] -6 * image_in[357] -24 * image_in[358] -38 * image_in[359] -1 * image_in[360] +26 * image_in[361] +4 * image_in[362] -11 * image_in[363] +2 * image_in[364] -19 * image_in[365] +6 * image_in[366] -24 * image_in[367] -83 * image_in[368] -101 * image_in[369] -82 * image_in[370] -67 * image_in[371] -19 * image_in[372] -12 * image_in[373] -26 * image_in[374] -31 * image_in[375] -25 * image_in[376] -5 * image_in[377] +3 * image_in[378] -10 * image_in[379] -5 * image_in[380] -2 * image_in[381] -6 * image_in[382] -6 * image_in[383]
                            -31 * image_in[384] -31 * image_in[385] -39 * image_in[386] -32 * image_in[387] -9 * image_in[388] +14 * image_in[389] +4 * image_in[390] +4 * image_in[391] +3 * image_in[392] +3 * image_in[393] +8 * image_in[394] -26 * image_in[395] -63 * image_in[396] -51 * image_in[397] -37 * image_in[398] -12 * image_in[399] -2 * image_in[400] -9 * image_in[401] -21 * image_in[402] -22 * image_in[403] +8 * image_in[405] +10 * image_in[406] +17 * image_in[407] -9 * image_in[408] -7 * image_in[409] -9 * image_in[410] -17 * image_in[411] -27 * image_in[412] -19 * image_in[413] -45 * image_in[414] -37 * image_in[415]
                            -20 * image_in[416] -13 * image_in[417] +29 * image_in[418] +3 * image_in[419] -1 * image_in[420] +16 * image_in[421] +26 * image_in[422] -22 * image_in[423] +2 * image_in[424] -6 * image_in[425] -11 * image_in[426] +5 * image_in[427] -6 * image_in[428] -7 * image_in[429] -8 * image_in[430] -12 * image_in[431] +4 * image_in[432] +12 * image_in[433] +15 * image_in[434] +8 * image_in[435] -6 * image_in[436] -14 * image_in[437] -17 * image_in[438] -21 * image_in[439] -19 * image_in[440] -19 * image_in[441] -18 * image_in[442] -16 * image_in[443] -6 * image_in[444] -11 * image_in[445] +19 * image_in[446] +7 * image_in[447]
                            -6 * image_in[448] -5 * image_in[449] +35 * image_in[450] +34 * image_in[451] +33 * image_in[452] +21 * image_in[453] -2 * image_in[454] -3 * image_in[455] -19 * image_in[456] +23 * image_in[457] +9 * image_in[458] +6 * image_in[459] +4 * image_in[460] +15 * image_in[461] -4 * image_in[462] -16 * image_in[463] -8 * image_in[464] -1 * image_in[465] -3 * image_in[466] -4 * image_in[467] -22 * image_in[468] -10 * image_in[469] -8 * image_in[470] +12 * image_in[472] +27 * image_in[473] +13 * image_in[474] +23 * image_in[475] +4 * image_in[476] +16 * image_in[477] +8 * image_in[478] +52 * image_in[479]
                            +44 * image_in[480] +11 * image_in[481] -5 * image_in[482] -11 * image_in[483] -1 * image_in[484] -4 * image_in[485] -5 * image_in[486] +1 * image_in[487] -17 * image_in[489] -32 * image_in[490] -22 * image_in[491] -3 * image_in[492] +2 * image_in[493] -5 * image_in[494] -3 * image_in[495] -22 * image_in[496] -24 * image_in[497] -9 * image_in[498] -14 * image_in[500] +22 * image_in[501] +50 * image_in[502] +1 * image_in[503] +1 * image_in[504] +13 * image_in[505] +41 * image_in[506] +25 * image_in[507] +17 * image_in[508] +7 * image_in[509] -5 * image_in[510] -8 * image_in[511]
                            -2 * image_in[512] +2 * image_in[513] +2 * image_in[514] -17 * image_in[515] -22 * image_in[516] -20 * image_in[517] -24 * image_in[518] -9 * image_in[519] +12 * image_in[520] +11 * image_in[521] +13 * image_in[522] +18 * image_in[523] -9 * image_in[524] -10 * image_in[525] +6 * image_in[526] +9 * image_in[527] +26 * image_in[528] +41 * image_in[529] +37 * image_in[530] +29 * image_in[531] +2 * image_in[532] +6 * image_in[533] -19 * image_in[534] +23 * image_in[535] +11 * image_in[536] +3 * image_in[537] -4 * image_in[538] -3 * image_in[539] +16 * image_in[540] +13 * image_in[541] +8 * image_in[542] -17 * image_in[543]
                            -9 * image_in[544] -11 * image_in[545] +4 * image_in[546] +2 * image_in[547] +11 * image_in[548] +20 * image_in[549] +9 * image_in[550] +1 * image_in[551] -3 * image_in[552] +10 * image_in[553] +3 * image_in[554] +6 * image_in[555] +4 * image_in[556] +37 * image_in[557] +28 * image_in[558] +19 * image_in[559] -1 * image_in[560] +20 * image_in[561] -4 * image_in[562] +23 * image_in[563] +20 * image_in[564] +20 * image_in[565] +22 * image_in[566] +19 * image_in[567] +17 * image_in[568] +22 * image_in[569] +25 * image_in[570] +4 * image_in[571] +3 * image_in[572] +5 * image_in[573] +14 * image_in[574] +12 * image_in[575]
                            +5 * image_in[576] +13 * image_in[577] +11 * image_in[578] +5 * image_in[579] +8 * image_in[580] +10 * image_in[581] -25 * image_in[582] -12 * image_in[583] +14 * image_in[584] +10 * image_in[585] -12 * image_in[586] +3 * image_in[587] +1 * image_in[588] +17 * image_in[589] +30 * image_in[590] +37 * image_in[591] +23 * image_in[592] +9 * image_in[593] +22 * image_in[594] +26 * image_in[595] +9 * image_in[596] +3 * image_in[597] +7 * image_in[598] +16 * image_in[599] +8 * image_in[600] +13 * image_in[601] +6 * image_in[602] +3 * image_in[603] +9 * image_in[604] +8 * image_in[605] +17 * image_in[606] +25 * image_in[607]
                            -8 * image_in[608] +4 * image_in[609] -10 * image_in[610] -11 * image_in[611] -2 * image_in[612] +22 * image_in[613] -25 * image_in[614] -1 * image_in[615] -3 * image_in[616] +1 * image_in[617] +34 * image_in[618] +41 * image_in[619] +11 * image_in[620] +10 * image_in[621] +30 * image_in[622] +22 * image_in[623] +4 * image_in[624] +15 * image_in[625] +9 * image_in[626] +17 * image_in[627] +14 * image_in[628] +17 * image_in[629] +5 * image_in[630] +19 * image_in[631] +11 * image_in[632] +8 * image_in[633] +11 * image_in[634] +24 * image_in[635] -7 * image_in[636] -7 * image_in[637] -3 * image_in[638] -4 * image_in[639]
                            +1 * image_in[640] -2 * image_in[641] +6 * image_in[642] -3 * image_in[643] -6 * image_in[644] +24 * image_in[646] +29 * image_in[647] +32 * image_in[648] +7 * image_in[649] +31 * image_in[650] +34 * image_in[651] +21 * image_in[652] +29 * image_in[653] +22 * image_in[654] +28 * image_in[655] +31 * image_in[656] +30 * image_in[657] +23 * image_in[658] +21 * image_in[659] +12 * image_in[660] +10 * image_in[661] +13 * image_in[662] -3 * image_in[663] -5 * image_in[664] -34 * image_in[665] +21 * image_in[667] +6 * image_in[668] -10 * image_in[669] -11 * image_in[670] -3 * image_in[671]
                            -2 * image_in[672] -3 * image_in[673] +20 * image_in[674] +28 * image_in[675] +41 * image_in[676] +20 * image_in[677] +18 * image_in[678] +25 * image_in[679] +12 * image_in[680] +8 * image_in[681] +20 * image_in[682] +29 * image_in[683] +30 * image_in[684] +44 * image_in[685] +32 * image_in[686] +19 * image_in[687] +27 * image_in[688] +25 * image_in[689] +1 * image_in[690] -16 * image_in[691] -37 * image_in[692] -18 * image_in[693] -20 * image_in[694] -23 * image_in[695] +14 * image_in[696] +22 * image_in[697] +4 * image_in[698] +3 * image_in[699] +5 * image_in[700] +2 * image_in[701] -4 * image_in[702] -18 * image_in[703]
                            +1 * image_in[704] +22 * image_in[706] +22 * image_in[707] +47 * image_in[708] +26 * image_in[709] +35 * image_in[710] +30 * image_in[711] +39 * image_in[712] +28 * image_in[713] +27 * image_in[714] +23 * image_in[715] +31 * image_in[716] +22 * image_in[717] +8 * image_in[718] +7 * image_in[719] -31 * image_in[720] -34 * image_in[721] -30 * image_in[722] -19 * image_in[723] -9 * image_in[724] +1 * image_in[725] -2 * image_in[726] +5 * image_in[727] +6 * image_in[728] -2 * image_in[729] +6 * image_in[730] +1 * image_in[731] -25 * image_in[732] -37 * image_in[733] -27 * image_in[734] +7 * image_in[735]
                            +14 * image_in[736] +4 * image_in[738] -4 * image_in[739] -21 * image_in[740] +4 * image_in[741] +22 * image_in[743] +34 * image_in[744] +24 * image_in[745] +14 * image_in[746] +20 * image_in[747] -9 * image_in[748] -17 * image_in[749] -10 * image_in[750] -1 * image_in[751] -5 * image_in[752] +1 * image_in[753] +1 * image_in[754] +1 * image_in[755] +4 * image_in[756] -1 * image_in[757] +1 * image_in[758] +3 * image_in[759] +4 * image_in[760] +20 * image_in[761] +24 * image_in[762] +27 * image_in[763] +26 * image_in[764] +2 * image_in[765] +15 * image_in[766] +3 * image_in[767] +31 * image_in[769] +17 * image_in[770] +36 * image_in[771] +18 * image_in[772] +37 * image_in[773] -6 * image_in[774] +11 * image_in[775] -5 * image_in[776] -23 * image_in[778] +1 * image_in[779] -5 * image_in[780] -1 * image_in[781] +4 * image_in[782] -3 * image_in[783];
                        if (layer1_out[1] < 0) layer1_out[1] = 0;
                        layer1_out[2] = 6 -5 * image_in[0] -2 * image_in[1] -1 * image_in[2] +6 * image_in[3] -4 * image_in[4] -1 * image_in[6] +6 * image_in[7] +2 * image_in[9] +5 * image_in[10] +4 * image_in[11] +4 * image_in[12] -15 * image_in[13] -3 * image_in[14] -4 * image_in[15] +2 * image_in[16] +2 * image_in[17] +4 * image_in[18] -1 * image_in[19] +3 * image_in[20] +4 * image_in[21] -1 * image_in[22] +6 * image_in[23] -1 * image_in[24] -3 * image_in[25] +4 * image_in[26] -4 * image_in[27] -5 * image_in[28] -5 * image_in[29] +5 * image_in[30] -6 * image_in[31]
                            -5 * image_in[32] -5 * image_in[33] -12 * image_in[34] -36 * image_in[35] -28 * image_in[36] -4 * image_in[37] -5 * image_in[38] -26 * image_in[39] -46 * image_in[40] -29 * image_in[41] -7 * image_in[42] -33 * image_in[43] -53 * image_in[44] -29 * image_in[45] -14 * image_in[47] -29 * image_in[48] -18 * image_in[49] -26 * image_in[50] -14 * image_in[51] -2 * image_in[52] +2 * image_in[53] +5 * image_in[54] -1 * image_in[55] +2 * image_in[56] -6 * image_in[57] -2 * image_in[58] -2 * image_in[59] -3 * image_in[61] -18 * image_in[62] -43 * image_in[63]
                            -36 * image_in[64] -31 * image_in[65] -54 * image_in[66] -25 * image_in[67] -47 * image_in[68] -16 * image_in[69] -15 * image_in[70] -27 * image_in[71] -42 * image_in[72] -38 * image_in[73] -29 * image_in[74] -3 * image_in[75] -7 * image_in[76] -25 * image_in[77] -17 * image_in[78] -32 * image_in[79] -20 * image_in[80] -16 * image_in[81] -2 * image_in[82] -3 * image_in[83] -6 * image_in[84] -3 * image_in[85] -14 * image_in[86] -1 * image_in[88] +11 * image_in[89] -14 * image_in[90] -16 * image_in[91] -25 * image_in[92] -40 * image_in[93] -24 * image_in[94] -18 * image_in[95]
                            -36 * image_in[96] -54 * image_in[97] -18 * image_in[98] -27 * image_in[99] -31 * image_in[100] -18 * image_in[101] +4 * image_in[102] -9 * image_in[103] -14 * image_in[104] +9 * image_in[105] +19 * image_in[106] +5 * image_in[107] -19 * image_in[108] +2 * image_in[110] -2 * image_in[111] +2 * image_in[112] -2 * image_in[113] -23 * image_in[114] +5 * image_in[115] +10 * image_in[116] +4 * image_in[117] -15 * image_in[118] -2 * image_in[119] -15 * image_in[120] -14 * image_in[121] -17 * image_in[122] -6 * image_in[123] -3 * image_in[124] -13 * image_in[125] -5 * image_in[126] +1 * image_in[127] -8 * image_in[129] -14 * image_in[130] +5 * image_in[131] +2 * image_in[132] +5 * image_in[133] +4 * image_in[134] +1 * image_in[135] +59 * image_in[136] +16 * image_in[137] +23 * image_in[138] -2 * image_in[139] -1 * image_in[140] -6 * image_in[141] -5 * image_in[142] -6 * image_in[143] -4 * image_in[144] +21 * image_in[145] +5 * image_in[146] +14 * image_in[147] +19 * image_in[148] +30 * image_in[149] -2 * image_in[150] +30 * image_in[151] +25 * image_in[152] +16 * image_in[153] +6 * image_in[154] +6 * image_in[155] -4 * image_in[156] -10 * image_in[157] -31 * image_in[158] -1 * image_in[159]
                            -17 * image_in[160] -29 * image_in[161] -33 * image_in[162] -11 * image_in[163] +5 * image_in[164] +22 * image_in[165] +7 * image_in[166] -5 * image_in[167] +3 * image_in[168] -3 * image_in[169] +30 * image_in[170] -4 * image_in[171] +16 * image_in[172] +1 * image_in[173] +1 * image_in[174] +7 * image_in[175] +30 * image_in[176] +21 * image_in[177] +26 * image_in[178] +30 * image_in[179] +26 * image_in[180] +17 * image_in[181] +19 * image_in[182] +27 * image_in[183] +7 * image_in[184] +18 * image_in[185] -5 * image_in[186] +5 * image_in[187] +4 * image_in[188] -15 * image_in[189] -9 * image_in[190] -10 * image_in[191]
                            -7 * image_in[192] +26 * image_in[193] +5 * image_in[194] -2 * image_in[195] -5 * image_in[196] -39 * image_in[197] +8 * image_in[198] +17 * image_in[199] -15 * image_in[200] -8 * image_in[201] +27 * image_in[203] +23 * image_in[204] +39 * image_in[205] +21 * image_in[206] +21 * image_in[207] +32 * image_in[208] +27 * image_in[209] +16 * image_in[210] +40 * image_in[211] +30 * image_in[212] +30 * image_in[213] +14 * image_in[214] +5 * image_in[215] +8 * image_in[216] -6 * image_in[217] -16 * image_in[218] +4 * image_in[219] +1 * image_in[220] +13 * image_in[221] -1 * image_in[222] +3 * image_in[223]
                            +13 * image_in[224] +18 * image_in[226] +6 * image_in[227] -4 * image_in[228] +17 * image_in[229] +23 * image_in[230] +28 * image_in[231] +37 * image_in[232] +29 * image_in[233] +11 * image_in[234] +22 * image_in[235] +15 * image_in[236] +17 * image_in[237] +4 * image_in[238] +8 * image_in[239] +9 * image_in[240] +1 * image_in[241] +21 * image_in[242] -6 * image_in[243] -4 * image_in[244] +10 * image_in[245] -7 * image_in[246] -15 * image_in[247] +23 * image_in[248] +17 * image_in[249] +3 * image_in[250] -6 * image_in[252] +6 * image_in[253] +19 * image_in[254] +5 * image_in[255]
                            -7 * image_in[256] +9 * image_in[257] +34 * image_in[258] +23 * image_in[259] +29 * image_in[260] +22 * image_in[261] +15 * image_in[262] +23 * image_in[263] +31 * image_in[264] +12 * image_in[265] -9 * image_in[266] -17 * image_in[267] -8 * image_in[268] -1 * image_in[269] -3 * image_in[270] +14 * image_in[271] +20 * image_in[272] +20 * image_in[273] +11 * image_in[274] -1 * image_in[275] -32 * image_in[276] -16 * image_in[277] +7 * image_in[278] +12 * image_in[279] +6 * image_in[280] +4 * image_in[281] -2 * image_in[282] -8 * image_in[283] +5 * image_in[284] +3 * image_in[285] +15 * image_in[286] +39 * image_in[287]
                            +40 * image_in[288] +38 * image_in[289] +42 * image_in[290] +33 * image_in[291] +25 * image_in[292] -2 * image_in[293] -30 * image_in[294] -35 * image_in[295] -20 * image_in[296] -18 * image_in[297] +6 * image_in[298] +25 * image_in[299] +21 * image_in[300] +18 * image_in[301] +20 * image_in[302] -15 * image_in[303] -62 * image_in[304] -46 * image_in[305] -30 * image_in[306] +16 * image_in[307] +1 * image_in[308] +8 * image_in[309] -17 * image_in[310] +24 * image_in[311] +18 * image_in[313] +30 * image_in[314] +50 * image_in[315] +42 * image_in[316] +66 * image_in[317] +79 * image_in[318] +58 * image_in[319]
                            +45 * image_in[320] -2 * image_in[321] +1 * image_in[322] +22 * image_in[323] +28 * image_in[324] +31 * image_in[325] +17 * image_in[326] +11 * image_in[327] +38 * image_in[328] +36 * image_in[329] +31 * image_in[330] -2 * image_in[331] -15 * image_in[332] -12 * image_in[333] +21 * image_in[334] +22 * image_in[335] +6 * image_in[336] +17 * image_in[337] +8 * image_in[338] +4 * image_in[339] +22 * image_in[340] +38 * image_in[341] +46 * image_in[342] +64 * image_in[343] +61 * image_in[344] +59 * image_in[345] +46 * image_in[346] +59 * image_in[347] +19 * image_in[348] +5 * image_in[349] +3 * image_in[350] +42 * image_in[351]
                            +55 * image_in[352] +46 * image_in[353] +32 * image_in[354] +24 * image_in[355] +43 * image_in[356] +52 * image_in[357] +49 * image_in[358] +37 * image_in[359] -6 * image_in[360] -18 * image_in[361] -27 * image_in[362] +16 * image_in[363] -3 * image_in[364] +13 * image_in[365] -17 * image_in[366] +7 * image_in[367] +44 * image_in[368] +48 * image_in[369] +44 * image_in[370] +71 * image_in[371] +37 * image_in[372] +38 * image_in[373] +37 * image_in[374] +21 * image_in[375] -11 * image_in[376] +4 * image_in[377] +7 * image_in[378] +56 * image_in[379] +63 * image_in[380] +39 * image_in[381] +35 * image_in[382] +23 * image_in[383]
                            +54 * image_in[384] +47 * image_in[385] +40 * image_in[386] +12 * image_in[387] -15 * image_in[388] -48 * image_in[389] -37 * image_in[390] -25 * image_in[391] +4 * image_in[392] +4 * image_in[393] +1 * image_in[394] +13 * image_in[395] +66 * image_in[396] +25 * image_in[397] +28 * image_in[398] +13 * image_in[399] +13 * image_in[400] +9 * image_in[401] +24 * image_in[402] +18 * image_in[403] +3 * image_in[404] +6 * image_in[405] +10 * image_in[406] +29 * image_in[407] +45 * image_in[408] +52 * image_in[409] +28 * image_in[410] +35 * image_in[411] +21 * image_in[412] +14 * image_in[413] +22 * image_in[414] -6 * image_in[415]
                            -50 * image_in[416] -35 * image_in[417] -39 * image_in[418] -4 * image_in[419] +1 * image_in[420] +17 * image_in[421] +6 * image_in[422] +11 * image_in[423] -9 * image_in[424] -17 * image_in[425] +4 * image_in[427] +4 * image_in[428] +5 * image_in[429] +15 * image_in[430] +7 * image_in[431] +17 * image_in[432] +13 * image_in[433] +6 * image_in[434] +34 * image_in[435] +37 * image_in[436] +40 * image_in[437] +24 * image_in[438] +11 * image_in[439] +18 * image_in[440] +9 * image_in[441] +22 * image_in[442] +2 * image_in[443] -67 * image_in[444] -57 * image_in[445] -39 * image_in[446] -15 * image_in[447]
                            +6 * image_in[448] +6 * image_in[449] +5 * image_in[450] -44 * image_in[451] -40 * image_in[452] -40 * image_in[453] -3 * image_in[454] +9 * image_in[455] +37 * image_in[456] +18 * image_in[457] +16 * image_in[458] +7 * image_in[459] +18 * image_in[460] +1 * image_in[461] -6 * image_in[462] +26 * image_in[463] +30 * image_in[464] +19 * image_in[465] +11 * image_in[466] +1 * image_in[468] -34 * image_in[469] -9 * image_in[470] -17 * image_in[471] -46 * image_in[472] -67 * image_in[473] -46 * image_in[474] -37 * image_in[475] -3 * image_in[476] +10 * image_in[477] -14 * image_in[478] -52 * image_in[479]
                            -51 * image_in[480] -51 * image_in[481] -33 * image_in[482] +2 * image_in[483] +21 * image_in[484] +30 * image_in[485] +4 * image_in[486] +6 * image_in[487] +13 * image_in[488] +5 * image_in[489] +10 * image_in[490] +11 * image_in[491] +28 * image_in[492] +18 * image_in[493] +8 * image_in[494] -1 * image_in[495] +4 * image_in[496] +10 * image_in[497] -5 * image_in[498] -14 * image_in[499] -34 * image_in[500] -70 * image_in[501] -53 * image_in[502] -5 * image_in[503] +4 * image_in[504] +8 * image_in[505] -12 * image_in[506] -37 * image_in[507] -47 * image_in[508] -46 * image_in[509] -25 * image_in[510] -20 * image_in[511]
                            -3 * image_in[512] +8 * image_in[513] -7 * image_in[514] -4 * image_in[515] -12 * image_in[516] -13 * image_in[517] -6 * image_in[518] +13 * image_in[519] +5 * image_in[520] -10 * image_in[521] +2 * image_in[522] +4 * image_in[523] +18 * image_in[524] +2 * image_in[525] -22 * image_in[526] -30 * image_in[527] -78 * image_in[528] -78 * image_in[529] -37 * image_in[530] -20 * image_in[531] -5 * image_in[532] +9 * image_in[533] -1 * image_in[534] -32 * image_in[535] -42 * image_in[536] -14 * image_in[537] -32 * image_in[538] -32 * image_in[539] -24 * image_in[540] -34 * image_in[541] -32 * image_in[542] -33 * image_in[543]
                            -31 * image_in[544] -40 * image_in[545] -15 * image_in[546] -15 * image_in[547] -8 * image_in[548] -4 * image_in[549] -7 * image_in[550] +22 * image_in[551] +7 * image_in[552] +2 * image_in[553] -23 * image_in[554] -13 * image_in[555] -19 * image_in[556] -67 * image_in[557] -32 * image_in[558] -5 * image_in[559] -2 * image_in[560] -12 * image_in[561] +8 * image_in[562] -35 * image_in[563] -32 * image_in[564] -35 * image_in[565] -35 * image_in[566] -40 * image_in[567] -42 * image_in[568] -40 * image_in[569] -38 * image_in[570] -36 * image_in[571] -37 * image_in[572] -14 * image_in[573] -5 * image_in[574] +8 * image_in[575]
                            +6 * image_in[576] +7 * image_in[577] -2 * image_in[578] +10 * image_in[579] +6 * image_in[580] -6 * image_in[581] -14 * image_in[582] -17 * image_in[583] -27 * image_in[584] -19 * image_in[585] -22 * image_in[586] +4 * image_in[587] -1 * image_in[588] -6 * image_in[589] -31 * image_in[590] -74 * image_in[591] -58 * image_in[592] -29 * image_in[593] -28 * image_in[594] -31 * image_in[595] -27 * image_in[596] -17 * image_in[597] -25 * image_in[598] -19 * image_in[599] -7 * image_in[600] -9 * image_in[601] +8 * image_in[603] +11 * image_in[604] +5 * image_in[605] -1 * image_in[607]
                            +5 * image_in[608] -7 * image_in[609] -20 * image_in[610] -38 * image_in[611] -15 * image_in[612] -36 * image_in[613] -12 * image_in[614] -5 * image_in[615] +5 * image_in[616] +6 * image_in[617] -38 * image_in[618] -45 * image_in[619] -23 * image_in[620] -37 * image_in[621] -42 * image_in[622] -17 * image_in[623] -17 * image_in[624] -17 * image_in[625] -4 * image_in[626] -1 * image_in[627] +23 * image_in[628] +27 * image_in[629] +12 * image_in[630] +20 * image_in[631] +9 * image_in[632] +7 * image_in[633] -7 * image_in[634] +3 * image_in[635] -23 * image_in[636] -11 * image_in[637] -21 * image_in[638] +9 * image_in[639]
                            +8 * image_in[640] -10 * image_in[641] -19 * image_in[642] +4 * image_in[643] +2 * image_in[644] -5 * image_in[645] -20 * image_in[646] +9 * image_in[647] -9 * image_in[648] -23 * image_in[649] -18 * image_in[650] -13 * image_in[651] -5 * image_in[652] -13 * image_in[653] -7 * image_in[654] +2 * image_in[655] +9 * image_in[656] +19 * image_in[657] +31 * image_in[658] +15 * image_in[659] +21 * image_in[660] +16 * image_in[661] +8 * image_in[662] -10 * image_in[664] +3 * image_in[665] -4 * image_in[666] -7 * image_in[667] -13 * image_in[668] -14 * image_in[669] -22 * image_in[670] -6 * image_in[671]
                            +1 * image_in[672] +4 * image_in[673] -16 * image_in[674] +30 * image_in[675] +30 * image_in[677] +2 * image_in[678] +24 * image_in[679] +31 * image_in[680] +7 * image_in[681] +30 * image_in[682] +30 * image_in[683] +16 * image_in[684] +15 * image_in[685] +19 * image_in[686] +27 * image_in[687] +43 * image_in[688] +10 * image_in[689] +16 * image_in[690] +16 * image_in[691] +25 * image_in[692] -1 * image_in[693] +13 * image_in[694] +31 * image_in[695] -22 * image_in[696] -34 * image_in[697] -5 * image_in[698] +2 * image_in[699] +6 * image_in[700] -3 * image_in[701] +3 * image_in[702] -3 * image_in[703]
                            +18 * image_in[704] +38 * image_in[705] +13 * image_in[706] +32 * image_in[707] +24 * image_in[708] +42 * image_in[709] +56 * image_in[710] +55 * image_in[711] +32 * image_in[712] +36 * image_in[713] +39 * image_in[714] +42 * image_in[715] +37 * image_in[716] +28 * image_in[717] +39 * image_in[718] +28 * image_in[719] +41 * image_in[720] +34 * image_in[721] +5 * image_in[722] +4 * image_in[723] -10 * image_in[724] -6 * image_in[725] -1 * image_in[726] -1 * image_in[727] +3 * image_in[728] -2 * image_in[729] +5 * image_in[730] +3 * image_in[731] +34 * image_in[732] +56 * image_in[733] +27 * image_in[734] +39 * image_in[735]
                            +54 * image_in[736] +44 * image_in[737] +43 * image_in[738] +31 * image_in[739] +28 * image_in[740] +53 * image_in[741] +61 * image_in[742] +24 * image_in[743] +44 * image_in[744] +44 * image_in[745] +46 * image_in[746] +29 * image_in[747] +34 * image_in[748] +35 * image_in[749] +12 * image_in[750] +27 * image_in[751] -2 * image_in[752] -5 * image_in[753] -4 * image_in[754] -4 * image_in[755] +4 * image_in[756] +2 * image_in[757] +2 * image_in[758] +2 * image_in[759] +2 * image_in[760] -18 * image_in[761] -29 * image_in[762] +16 * image_in[763] +17 * image_in[764] +8 * image_in[765] +31 * image_in[766] -4 * image_in[767]
                            +4 * image_in[768] +42 * image_in[770] +35 * image_in[771] +28 * image_in[772] +17 * image_in[773] +32 * image_in[774] +17 * image_in[775] +18 * image_in[776] +23 * image_in[777] +29 * image_in[778] +1 * image_in[779] +2 * image_in[780] -2 * image_in[781] -1 * image_in[782] -2 * image_in[783];
                        if (layer1_out[2] < 0) layer1_out[2] = 0;
                        layer1_out[3] = -19 +2 * image_in[0] +5 * image_in[2] -3 * image_in[3] -1 * image_in[4] +1 * image_in[5] -1 * image_in[6] -5 * image_in[7] +6 * image_in[8] +1 * image_in[9] +4 * image_in[10] +4 * image_in[11] +2 * image_in[12] +7 * image_in[13] +9 * image_in[14] +4 * image_in[15] +4 * image_in[16] +1 * image_in[17] +1 * image_in[18] +4 * image_in[19] +2 * image_in[20] +1 * image_in[21] -1 * image_in[22] +3 * image_in[23] +2 * image_in[24] -2 * image_in[25] +6 * image_in[26] -3 * image_in[27] -6 * image_in[28] +5 * image_in[29] -5 * image_in[30] +5 * image_in[31]
                            -2 * image_in[32] +3 * image_in[33] -11 * image_in[34] -22 * image_in[35] -17 * image_in[36] -24 * image_in[37] -25 * image_in[38] -11 * image_in[39] -25 * image_in[40] -45 * image_in[41] +14 * image_in[42] +3 * image_in[43] +29 * image_in[44] -19 * image_in[45] -36 * image_in[46] -30 * image_in[47] -20 * image_in[48] -24 * image_in[49] -21 * image_in[50] -12 * image_in[51] -2 * image_in[52] +4 * image_in[53] +5 * image_in[54] -6 * image_in[55] -6 * image_in[56] -4 * image_in[57] +1 * image_in[58] -2 * image_in[59] -14 * image_in[60] -6 * image_in[61] -30 * image_in[62] -33 * image_in[63]
                            -29 * image_in[64] -14 * image_in[65] -36 * image_in[66] -18 * image_in[67] -28 * image_in[68] -48 * image_in[69] -72 * image_in[70] -60 * image_in[71] -58 * image_in[72] -48 * image_in[73] -44 * image_in[74] -46 * image_in[75] -43 * image_in[76] -45 * image_in[77] -33 * image_in[78] -21 * image_in[79] +11 * image_in[80] +16 * image_in[81] +6 * image_in[82] -6 * image_in[83] -4 * image_in[84] -3 * image_in[85] -13 * image_in[86] -1 * image_in[87] +1 * image_in[88] -12 * image_in[89] -38 * image_in[90] -26 * image_in[91] -10 * image_in[92] -7 * image_in[93] -18 * image_in[94] -14 * image_in[95]
                            -28 * image_in[96] -47 * image_in[97] -46 * image_in[98] -70 * image_in[99] -61 * image_in[100] -48 * image_in[101] -67 * image_in[102] -84 * image_in[103] -67 * image_in[104] -58 * image_in[105] -49 * image_in[106] -13 * image_in[107] +11 * image_in[108] +12 * image_in[109] +4 * image_in[110] -4 * image_in[111] +6 * image_in[112] +2 * image_in[113] +3 * image_in[114] +6 * image_in[115] -34 * image_in[116] -37 * image_in[117] -12 * image_in[118] -22 * image_in[119] -10 * image_in[120] -3 * image_in[122] -15 * image_in[123] +6 * image_in[124] -16 * image_in[125] -14 * image_in[126] -21 * image_in[127]
                            -38 * image_in[128] -31 * image_in[129] -18 * image_in[130] -23 * image_in[131] -19 * image_in[132] -33 * image_in[133] -42 * image_in[134] -24 * image_in[135] -20 * image_in[136] +2 * image_in[137] -11 * image_in[138] -5 * image_in[139] -1 * image_in[141] +4 * image_in[142] +22 * image_in[143] -7 * image_in[144] -23 * image_in[145] -29 * image_in[146] -16 * image_in[147] +2 * image_in[148] -6 * image_in[149] -8 * image_in[150] +36 * image_in[151] +24 * image_in[152] +31 * image_in[153] +11 * image_in[154] +5 * image_in[155] +3 * image_in[156] +9 * image_in[157] -8 * image_in[158] -14 * image_in[159]
                            -16 * image_in[160] -14 * image_in[161] -31 * image_in[162] -48 * image_in[163] -36 * image_in[164] +4 * image_in[165] -4 * image_in[166] -5 * image_in[168] +3 * image_in[169] +5 * image_in[170] +23 * image_in[171] -6 * image_in[172] -15 * image_in[173] -17 * image_in[174] -6 * image_in[175] +8 * image_in[176] +11 * image_in[177] +25 * image_in[178] +37 * image_in[179] +41 * image_in[180] +48 * image_in[181] +59 * image_in[182] +57 * image_in[183] +39 * image_in[184] +47 * image_in[185] +36 * image_in[186] +14 * image_in[187] +8 * image_in[188] +1 * image_in[189] -14 * image_in[190] -36 * image_in[191]
                            -59 * image_in[192] -7 * image_in[193] -21 * image_in[194] +6 * image_in[195] -3 * image_in[196] -37 * image_in[197] +38 * image_in[198] +36 * image_in[199] -7 * image_in[200] -31 * image_in[201] +2 * image_in[202] -10 * image_in[203] +3 * image_in[204] +23 * image_in[205] +21 * image_in[206] +33 * image_in[207] +45 * image_in[208] +51 * image_in[209] +47 * image_in[210] +58 * image_in[211] +51 * image_in[212] +34 * image_in[213] +28 * image_in[214] +13 * image_in[215] +9 * image_in[216] +4 * image_in[217] -2 * image_in[218] -14 * image_in[219] -9 * image_in[220] -30 * image_in[221] -26 * image_in[222] +10 * image_in[223]
                            +7 * image_in[224] +7 * image_in[225] -6 * image_in[226] +8 * image_in[227] +1 * image_in[228] -16 * image_in[229] +13 * image_in[230] +6 * image_in[231] +22 * image_in[232] +15 * image_in[233] +30 * image_in[234] +33 * image_in[235] +29 * image_in[236] +40 * image_in[237] +47 * image_in[238] +34 * image_in[239] +38 * image_in[240] +7 * image_in[241] +25 * image_in[242] +12 * image_in[243] +6 * image_in[244] +15 * image_in[245] +11 * image_in[246] +12 * image_in[247] -27 * image_in[249] -9 * image_in[250] -11 * image_in[251] +5 * image_in[252] +3 * image_in[253] -19 * image_in[254] +22 * image_in[255]
                            +2 * image_in[256] +21 * image_in[257] +27 * image_in[258] +2 * image_in[259] +9 * image_in[260] +31 * image_in[261] +33 * image_in[262] +22 * image_in[263] +41 * image_in[264] +46 * image_in[265] +27 * image_in[266] +16 * image_in[267] +25 * image_in[268] +23 * image_in[269] +29 * image_in[270] +28 * image_in[271] +23 * image_in[272] -3 * image_in[273] +3 * image_in[274] +18 * image_in[275] +3 * image_in[276] -26 * image_in[277] -6 * image_in[278] +21 * image_in[279] +8 * image_in[280] +5 * image_in[281] +17 * image_in[282] +7 * image_in[283] +14 * image_in[284] +29 * image_in[285] +45 * image_in[286] +14 * image_in[287]
                            +18 * image_in[288] +32 * image_in[289] +35 * image_in[290] +24 * image_in[291] +27 * image_in[292] +4 * image_in[293] +7 * image_in[294] -10 * image_in[295] -7 * image_in[296] +5 * image_in[297] +28 * image_in[298] +28 * image_in[299] +21 * image_in[300] +6 * image_in[301] +27 * image_in[302] +24 * image_in[303] -20 * image_in[304] -69 * image_in[305] -28 * image_in[306] +10 * image_in[307] +3 * image_in[308] +12 * image_in[309] +19 * image_in[310] +18 * image_in[311] +10 * image_in[312] +18 * image_in[313] +21 * image_in[314] +27 * image_in[315] +32 * image_in[316] +23 * image_in[317] +17 * image_in[318] +17 * image_in[319]
                            -12 * image_in[320] -9 * image_in[321] -10 * image_in[322] -28 * image_in[323] -13 * image_in[324] +18 * image_in[325] +24 * image_in[326] +21 * image_in[327] +36 * image_in[328] +30 * image_in[329] +38 * image_in[330] +19 * image_in[331] -9 * image_in[332] -18 * image_in[333] -4 * image_in[334] -21 * image_in[335] +7 * image_in[336] +18 * image_in[337] +21 * image_in[338] +17 * image_in[339] +24 * image_in[340] +26 * image_in[341] +4 * image_in[342] -1 * image_in[343] +11 * image_in[344] +5 * image_in[345] -11 * image_in[346] -17 * image_in[347] -42 * image_in[348] -29 * image_in[349] -18 * image_in[350] -32 * image_in[351]
                            -17 * image_in[352] +15 * image_in[353] +28 * image_in[354] +36 * image_in[355] +43 * image_in[356] +29 * image_in[357] +48 * image_in[358] +22 * image_in[359] +33 * image_in[360] +28 * image_in[361] +38 * image_in[362] -13 * image_in[363] +1 * image_in[364] +6 * image_in[365] +29 * image_in[366] +42 * image_in[367] +12 * image_in[368] -8 * image_in[369] -13 * image_in[370] -5 * image_in[371] -7 * image_in[373] -4 * image_in[374] -16 * image_in[375] -37 * image_in[376] -30 * image_in[377] -21 * image_in[378] -15 * image_in[379] +13 * image_in[380] +16 * image_in[381] +20 * image_in[382] +15 * image_in[383]
                            +21 * image_in[384] +18 * image_in[385] +20 * image_in[386] +16 * image_in[387] +24 * image_in[388] +43 * image_in[389] +37 * image_in[390] +25 * image_in[391] -2 * image_in[392] +17 * image_in[393] +4 * image_in[394] +17 * image_in[395] -15 * image_in[397] -9 * image_in[398] +15 * image_in[399] -7 * image_in[400] -12 * image_in[401] -7 * image_in[402] -5 * image_in[403] -28 * image_in[404] -2 * image_in[405] -25 * image_in[406] -9 * image_in[407] -6 * image_in[408] +22 * image_in[409] +23 * image_in[410] +14 * image_in[411] +8 * image_in[412] +10 * image_in[413] +4 * image_in[414] +8 * image_in[415]
                            +8 * image_in[416] +36 * image_in[417] +58 * image_in[418] +2 * image_in[419] -6 * image_in[420] -20 * image_in[421] -34 * image_in[422] +13 * image_in[423] +15 * image_in[424] +3 * image_in[425] -9 * image_in[428] -7 * image_in[429] -7 * image_in[430] -15 * image_in[431] -22 * image_in[432] -13 * image_in[433] -22 * image_in[434] +8 * image_in[436] +23 * image_in[437] +11 * image_in[438] +3 * image_in[440] -9 * image_in[441] +1 * image_in[442] -14 * image_in[443] +19 * image_in[444] +17 * image_in[445] +40 * image_in[446] +17 * image_in[447]
                            -5 * image_in[448] +1 * image_in[449] -24 * image_in[450] +4 * image_in[451] +20 * image_in[452] +1 * image_in[453] +12 * image_in[454] +17 * image_in[455] +5 * image_in[456] +1 * image_in[457] +6 * image_in[458] -4 * image_in[459] +7 * image_in[460] -13 * image_in[461] -12 * image_in[462] +1 * image_in[463] +27 * image_in[464] +35 * image_in[465] -25 * image_in[467] -5 * image_in[468] -3 * image_in[469] -4 * image_in[470] -10 * image_in[471] -14 * image_in[472] +38 * image_in[473] +60 * image_in[474] +37 * image_in[475] +6 * image_in[476] -10 * image_in[477] -28 * image_in[478] -10 * image_in[479]
                            +4 * image_in[480] -8 * image_in[481] +4 * image_in[482] +3 * image_in[483] +4 * image_in[484] +15 * image_in[485] +16 * image_in[486] +23 * image_in[487] +14 * image_in[488] -13 * image_in[490] +16 * image_in[491] +13 * image_in[492] +8 * image_in[493] -5 * image_in[494] -15 * image_in[495] -12 * image_in[496] -13 * image_in[497] -6 * image_in[498] -13 * image_in[499] +13 * image_in[500] +63 * image_in[501] +59 * image_in[502] +4 * image_in[503] -3 * image_in[505] -28 * image_in[506] -44 * image_in[507] -1 * image_in[508] -4 * image_in[509] +1 * image_in[510] +11 * image_in[511]
                            +2 * image_in[512] +10 * image_in[513] +32 * image_in[514] +20 * image_in[515] -17 * image_in[516] -15 * image_in[517] -10 * image_in[518] -2 * image_in[519] -7 * image_in[520] -9 * image_in[521] +4 * image_in[522] -14 * image_in[523] -12 * image_in[524] -16 * image_in[525] -12 * image_in[526] -7 * image_in[527] +25 * image_in[528] +30 * image_in[529] +11 * image_in[530] +37 * image_in[531] +3 * image_in[532] -45 * image_in[534] -46 * image_in[535] -14 * image_in[536] -7 * image_in[537] -5 * image_in[538] +15 * image_in[539] +11 * image_in[540] +2 * image_in[541] +6 * image_in[542] -20 * image_in[543]
                            -20 * image_in[544] -5 * image_in[545] -4 * image_in[546] -19 * image_in[547] -20 * image_in[548] -7 * image_in[549] -14 * image_in[550] -1 * image_in[551] -5 * image_in[552] -14 * image_in[553] +8 * image_in[554] +13 * image_in[555] -8 * image_in[556] +22 * image_in[557] +26 * image_in[558] +10 * image_in[559] -2 * image_in[560] +17 * image_in[561] -36 * image_in[562] -32 * image_in[563] -19 * image_in[564] +9 * image_in[565] -4 * image_in[566] +4 * image_in[567] +7 * image_in[568] -18 * image_in[569] -11 * image_in[570] -23 * image_in[571] -7 * image_in[572] -5 * image_in[573] -19 * image_in[574] -14 * image_in[575]
                            -16 * image_in[576] -26 * image_in[577] -23 * image_in[578] -13 * image_in[579] -22 * image_in[580] -12 * image_in[581] -4 * image_in[582] -6 * image_in[583] +20 * image_in[584] +9 * image_in[585] -9 * image_in[586] +5 * image_in[587] -5 * image_in[588] +1 * image_in[589] +11 * image_in[590] -26 * image_in[591] -10 * image_in[592] -4 * image_in[593] +5 * image_in[594] -9 * image_in[595] -8 * image_in[596] +3 * image_in[597] -6 * image_in[598] -2 * image_in[599] -3 * image_in[600] -20 * image_in[601] -15 * image_in[602] -19 * image_in[603] -9 * image_in[604] -26 * image_in[605] -22 * image_in[606] -20 * image_in[607]
                            -17 * image_in[608] -14 * image_in[609] -10 * image_in[610] +13 * image_in[611] +19 * image_in[612] +13 * image_in[613] -6 * image_in[614] +4 * image_in[615] +1 * image_in[616] -1 * image_in[617] -12 * image_in[618] -12 * image_in[619] -24 * image_in[620] -25 * image_in[621] +11 * image_in[622] +18 * image_in[623] +27 * image_in[624] +21 * image_in[625] +18 * image_in[626] +8 * image_in[627] +13 * image_in[628] +13 * image_in[629] -1 * image_in[630] -10 * image_in[631] +4 * image_in[632] -14 * image_in[633] -16 * image_in[634] -6 * image_in[635] -4 * image_in[637] +22 * image_in[638] +25 * image_in[639]
                            +29 * image_in[640] -3 * image_in[641] -11 * image_in[642] -6 * image_in[643] -2 * image_in[644] -4 * image_in[645] -21 * image_in[646] -23 * image_in[647] -32 * image_in[648] -23 * image_in[649] -16 * image_in[650] +12 * image_in[651] +25 * image_in[652] +9 * image_in[653] +21 * image_in[654] +16 * image_in[655] +21 * image_in[656] +16 * image_in[657] +13 * image_in[658] -1 * image_in[659] +4 * image_in[660] +9 * image_in[661] +1 * image_in[662] -4 * image_in[663] -3 * image_in[664] +36 * image_in[665] +47 * image_in[666] +33 * image_in[667] +29 * image_in[668] -4 * image_in[669] -14 * image_in[670] -5 * image_in[671]
                            -5 * image_in[672] -5 * image_in[673] -19 * image_in[674] -19 * image_in[675] -16 * image_in[676] +12 * image_in[677] -11 * image_in[678] +3 * image_in[679] +3 * image_in[680] -11 * image_in[681] +10 * image_in[682] -2 * image_in[683] +7 * image_in[684] +6 * image_in[685] +16 * image_in[687] +22 * image_in[688] +12 * image_in[689] +22 * image_in[690] +18 * image_in[691] +38 * image_in[692] +27 * image_in[693] +17 * image_in[694] +12 * image_in[695] +12 * image_in[696] +13 * image_in[697] +4 * image_in[698] +3 * image_in[699] +4 * image_in[700] -6 * image_in[701] +2 * image_in[702] -17 * image_in[703]
                            +9 * image_in[704] +17 * image_in[705] -6 * image_in[706] +23 * image_in[707] +1 * image_in[708] -2 * image_in[709] +8 * image_in[710] +20 * image_in[711] +6 * image_in[712] +16 * image_in[713] +14 * image_in[714] +28 * image_in[715] +32 * image_in[716] +29 * image_in[717] +26 * image_in[718] +32 * image_in[719] +43 * image_in[720] +38 * image_in[721] -11 * image_in[722] -5 * image_in[723] -10 * image_in[724] -2 * image_in[725] +5 * image_in[726] +2 * image_in[727] +5 * image_in[728] -6 * image_in[729] +4 * image_in[730] -5 * image_in[731] +30 * image_in[732] +28 * image_in[733] +24 * image_in[734] +49 * image_in[735]
                            +65 * image_in[736] +53 * image_in[737] +54 * image_in[738] +47 * image_in[739] +37 * image_in[740] +66 * image_in[741] +75 * image_in[742] +39 * image_in[743] +61 * image_in[744] +48 * image_in[745] +57 * image_in[746] +47 * image_in[747] +37 * image_in[748] +53 * image_in[749] +20 * image_in[750] +19 * image_in[751] +2 * image_in[752] -3 * image_in[753] -5 * image_in[754] +1 * image_in[755] -3 * image_in[756] -4 * image_in[757] -3 * image_in[758] +4 * image_in[759] +4 * image_in[760] -18 * image_in[761] -24 * image_in[762] +14 * image_in[763] +25 * image_in[764] +29 * image_in[765] +41 * image_in[766] +6 * image_in[767]
                            +17 * image_in[768] +6 * image_in[769] +52 * image_in[770] +44 * image_in[771] +37 * image_in[772] +18 * image_in[773] +38 * image_in[774] +30 * image_in[775] +17 * image_in[776] +27 * image_in[777] +24 * image_in[778] +5 * image_in[779] +4 * image_in[780] +6 * image_in[781] -2 * image_in[782] -1 * image_in[783];
                        if (layer1_out[3] < 0) layer1_out[3] = 0;
                        layer1_out[4] = 96 -1 * image_in[0] +4 * image_in[1] +1 * image_in[2] +2 * image_in[3] -2 * image_in[4] -3 * image_in[6] +4 * image_in[7] +3 * image_in[8] +6 * image_in[10] +3 * image_in[11] +3 * image_in[12] -14 * image_in[13] +1 * image_in[14] +4 * image_in[15] -1 * image_in[16] -1 * image_in[17] -2 * image_in[18] -3 * image_in[19] -4 * image_in[20] +2 * image_in[21] -2 * image_in[22] +5 * image_in[24] +5 * image_in[25] +1 * image_in[26] +3 * image_in[27] -5 * image_in[28] +4 * image_in[29] -5 * image_in[30] +3 * image_in[31]
                            -5 * image_in[32] -4 * image_in[34] -17 * image_in[35] -18 * image_in[36] +3 * image_in[38] -17 * image_in[39] -22 * image_in[40] -8 * image_in[41] +20 * image_in[42] +18 * image_in[43] -28 * image_in[44] +6 * image_in[45] +14 * image_in[46] -3 * image_in[47] -2 * image_in[48] -22 * image_in[49] -21 * image_in[50] -16 * image_in[51] +5 * image_in[52] -6 * image_in[53] -3 * image_in[54] -4 * image_in[55] -4 * image_in[56] +4 * image_in[57] +2 * image_in[58] +1 * image_in[59] -4 * image_in[60] -1 * image_in[61] +18 * image_in[62] -9 * image_in[63]
                            -5 * image_in[64] +10 * image_in[65] +31 * image_in[67] +27 * image_in[68] +71 * image_in[69] +68 * image_in[70] +55 * image_in[71] +38 * image_in[72] +29 * image_in[73] +1 * image_in[74] +12 * image_in[75] +33 * image_in[76] +17 * image_in[77] +25 * image_in[78] +19 * image_in[79] +20 * image_in[80] +12 * image_in[81] -3 * image_in[82] -2 * image_in[83] +1 * image_in[84] -2 * image_in[85] -12 * image_in[86] -1 * image_in[87] +23 * image_in[89] +33 * image_in[90] +44 * image_in[91] +23 * image_in[92] +9 * image_in[93] +40 * image_in[94] +32 * image_in[95]
                            +29 * image_in[96] +27 * image_in[97] +14 * image_in[98] +21 * image_in[99] +17 * image_in[100] +16 * image_in[101] +17 * image_in[102] +37 * image_in[103] +16 * image_in[104] -2 * image_in[105] -9 * image_in[106] -8 * image_in[107] +7 * image_in[108] -22 * image_in[109] +6 * image_in[110] -5 * image_in[111] -5 * image_in[112] +2 * image_in[113] +22 * image_in[114] -4 * image_in[115] +26 * image_in[116] +71 * image_in[117] +54 * image_in[118] +36 * image_in[119] +36 * image_in[120] +26 * image_in[121] +24 * image_in[122] +18 * image_in[123] +17 * image_in[124] +20 * image_in[125] +6 * image_in[126] -13 * image_in[127]
                            +1 * image_in[128] -5 * image_in[129] +10 * image_in[131] +20 * image_in[132] -9 * image_in[133] +15 * image_in[134] -8 * image_in[135] -28 * image_in[136] -22 * image_in[137] -17 * image_in[138] -5 * image_in[139] -4 * image_in[140] +3 * image_in[141] +5 * image_in[142] +12 * image_in[143] +50 * image_in[144] +54 * image_in[145] +50 * image_in[146] +23 * image_in[147] +6 * image_in[148] +14 * image_in[149] +13 * image_in[150] +9 * image_in[151] +19 * image_in[152] +13 * image_in[153] +10 * image_in[154] +11 * image_in[155] +13 * image_in[156] -2 * image_in[157] +12 * image_in[158] +12 * image_in[159]
                            -2 * image_in[160] +1 * image_in[161] +13 * image_in[162] +24 * image_in[163] -2 * image_in[164] -35 * image_in[165] +2 * image_in[166] -5 * image_in[167] +2 * image_in[168] -2 * image_in[169] -12 * image_in[170] +14 * image_in[171] +25 * image_in[172] +22 * image_in[173] +24 * image_in[174] +8 * image_in[175] +1 * image_in[176] +20 * image_in[177] +22 * image_in[178] +17 * image_in[179] +9 * image_in[180] +16 * image_in[181] +26 * image_in[182] -2 * image_in[183] +9 * image_in[184] -3 * image_in[185] +19 * image_in[186] -4 * image_in[187] -8 * image_in[188] -13 * image_in[189] -8 * image_in[190] +2 * image_in[191]
                            -26 * image_in[192] -49 * image_in[193] +5 * image_in[194] -4 * image_in[196] +28 * image_in[197] -27 * image_in[198] +36 * image_in[200] +9 * image_in[201] +15 * image_in[202] -10 * image_in[203] -9 * image_in[204] +13 * image_in[206] +8 * image_in[207] +19 * image_in[208] +27 * image_in[209] +41 * image_in[210] +13 * image_in[211] +4 * image_in[212] -11 * image_in[214] +2 * image_in[215] -11 * image_in[217] -17 * image_in[218] -54 * image_in[219] -67 * image_in[220] -29 * image_in[221] +11 * image_in[222] -14 * image_in[223]
                            -7 * image_in[224] -17 * image_in[225] -10 * image_in[226] -5 * image_in[227] +24 * image_in[228] -2 * image_in[229] -22 * image_in[230] -24 * image_in[231] -14 * image_in[232] -12 * image_in[233] -1 * image_in[234] +10 * image_in[235] -11 * image_in[236] +9 * image_in[237] +19 * image_in[238] +14 * image_in[239] -11 * image_in[240] +2 * image_in[241] -16 * image_in[242] -6 * image_in[243] -22 * image_in[244] -21 * image_in[245] -35 * image_in[246] -82 * image_in[247] -100 * image_in[248] -48 * image_in[249] -49 * image_in[250] -27 * image_in[251] -11 * image_in[252] -10 * image_in[253] -12 * image_in[254] -14 * image_in[255]
                            +4 * image_in[256] -24 * image_in[257] -28 * image_in[258] -11 * image_in[259] -18 * image_in[260] -2 * image_in[261] -5 * image_in[262] -6 * image_in[263] -7 * image_in[264] -5 * image_in[265] +2 * image_in[266] +40 * image_in[267] +7 * image_in[268] +1 * image_in[269] -10 * image_in[270] -18 * image_in[271] -25 * image_in[272] -29 * image_in[273] -29 * image_in[274] -59 * image_in[275] -91 * image_in[276] -84 * image_in[277] -42 * image_in[278] +14 * image_in[279] -16 * image_in[280] -17 * image_in[281] -33 * image_in[282] -4 * image_in[283] -42 * image_in[284] -14 * image_in[285] -18 * image_in[286] -11 * image_in[287]
                            -8 * image_in[288] -23 * image_in[289] -22 * image_in[290] -21 * image_in[291] -22 * image_in[292] -27 * image_in[293] -19 * image_in[294] +23 * image_in[295] +22 * image_in[296] +20 * image_in[297] -9 * image_in[298] -13 * image_in[299] -29 * image_in[300] -38 * image_in[301] -40 * image_in[302] -71 * image_in[303] -92 * image_in[304] -57 * image_in[305] -51 * image_in[306] -15 * image_in[307] -8 * image_in[308] -29 * image_in[309] -50 * image_in[310] -6 * image_in[311] -32 * image_in[312] -11 * image_in[313] -32 * image_in[314] -42 * image_in[315] -23 * image_in[316] -12 * image_in[317] -9 * image_in[318] -13 * image_in[319]
                            -27 * image_in[320] -39 * image_in[321] -24 * image_in[322] +15 * image_in[323] +32 * image_in[324] +26 * image_in[325] +9 * image_in[326] +8 * image_in[327] -1 * image_in[328] -24 * image_in[329] -44 * image_in[330] -64 * image_in[331] -73 * image_in[332] -62 * image_in[333] -55 * image_in[334] +14 * image_in[335] -8 * image_in[336] -25 * image_in[337] -40 * image_in[338] -42 * image_in[339] -29 * image_in[340] -12 * image_in[341] -13 * image_in[342] -12 * image_in[343] -6 * image_in[344] +1 * image_in[345] +3 * image_in[346] -5 * image_in[347] -4 * image_in[348] -7 * image_in[349] +21 * image_in[350] +31 * image_in[351]
                            +47 * image_in[352] +24 * image_in[353] +9 * image_in[354] +10 * image_in[355] -11 * image_in[356] -15 * image_in[357] -23 * image_in[358] -17 * image_in[359] -20 * image_in[360] -28 * image_in[361] -50 * image_in[362] +19 * image_in[363] +1 * image_in[364] -8 * image_in[365] -45 * image_in[366] -39 * image_in[367] -4 * image_in[369] +7 * image_in[370] -6 * image_in[371] +20 * image_in[372] +12 * image_in[373] +1 * image_in[375] +16 * image_in[376] +29 * image_in[377] +50 * image_in[378] +46 * image_in[379] +46 * image_in[380] +42 * image_in[381] +17 * image_in[382] +5 * image_in[383]
                            -5 * image_in[384] +1 * image_in[385] -10 * image_in[386] -9 * image_in[388] -9 * image_in[389] -5 * image_in[390] +12 * image_in[391] +1 * image_in[392] -13 * image_in[393] -29 * image_in[394] +5 * image_in[395] +16 * image_in[396] +15 * image_in[397] +14 * image_in[398] +20 * image_in[399] +28 * image_in[400] +19 * image_in[401] -3 * image_in[402] +18 * image_in[403] +30 * image_in[404] +32 * image_in[405] +50 * image_in[406] +53 * image_in[407] +58 * image_in[408] +33 * image_in[409] +18 * image_in[410] +3 * image_in[411] +11 * image_in[412] -3 * image_in[414] +3 * image_in[415]
                            -12 * image_in[416] +15 * image_in[417] +12 * image_in[418] +3 * image_in[419] +1 * image_in[420] +11 * image_in[421] -17 * image_in[422] +12 * image_in[423] +18 * image_in[424] +29 * image_in[425] +41 * image_in[426] +17 * image_in[427] +21 * image_in[428] +1 * image_in[429] +2 * image_in[430] +26 * image_in[431] +37 * image_in[432] +41 * image_in[433] +61 * image_in[434] +56 * image_in[435] +60 * image_in[436] +26 * image_in[437] -9 * image_in[438] +11 * image_in[439] -6 * image_in[440] +4 * image_in[441] +12 * image_in[442] -4 * image_in[443] -22 * image_in[444] +11 * image_in[445] +36 * image_in[446] +18 * image_in[447]
                            +4 * image_in[448] -2 * image_in[449] +48 * image_in[450] +8 * image_in[451] +13 * image_in[452] +51 * image_in[453] +25 * image_in[454] +16 * image_in[455] -6 * image_in[456] +10 * image_in[458] +20 * image_in[459] +28 * image_in[460] +53 * image_in[461] +63 * image_in[462] +36 * image_in[463] +38 * image_in[464] +11 * image_in[465] +14 * image_in[466] +13 * image_in[467] +11 * image_in[468] +15 * image_in[469] +21 * image_in[470] +4 * image_in[471] +31 * image_in[472] +42 * image_in[473] +48 * image_in[474] +28 * image_in[475] +1 * image_in[476] +16 * image_in[477] +52 * image_in[478] +36 * image_in[479]
                            +14 * image_in[480] +8 * image_in[481] -14 * image_in[482] +2 * image_in[483] -7 * image_in[484] -31 * image_in[485] -13 * image_in[486] -13 * image_in[487] +21 * image_in[488] +39 * image_in[489] +44 * image_in[490] +36 * image_in[491] +10 * image_in[492] +4 * image_in[493] +8 * image_in[494] +15 * image_in[495] +16 * image_in[496] +28 * image_in[497] +13 * image_in[498] +19 * image_in[499] -37 * image_in[500] +43 * image_in[501] +43 * image_in[502] +4 * image_in[503] -5 * image_in[504] +6 * image_in[505] +36 * image_in[506] +50 * image_in[507] +16 * image_in[508] +6 * image_in[509] -7 * image_in[510] -18 * image_in[511]
                            -36 * image_in[512] -39 * image_in[513] -37 * image_in[514] -20 * image_in[515] +17 * image_in[516] +17 * image_in[517] +37 * image_in[518] +23 * image_in[519] +30 * image_in[520] +26 * image_in[521] +27 * image_in[522] +19 * image_in[523] +25 * image_in[524] +27 * image_in[525] -2 * image_in[526] +7 * image_in[527] +13 * image_in[528] +65 * image_in[529] +47 * image_in[530] +24 * image_in[531] -2 * image_in[532] +13 * image_in[533] +1 * image_in[534] +53 * image_in[535] +14 * image_in[536] -11 * image_in[537] -13 * image_in[538] -5 * image_in[539] -33 * image_in[540] -36 * image_in[541] -37 * image_in[542] -3 * image_in[543]
                            -18 * image_in[544] +14 * image_in[545] +20 * image_in[546] +33 * image_in[547] +42 * image_in[548] +36 * image_in[549] +35 * image_in[550] +28 * image_in[551] +12 * image_in[552] +28 * image_in[553] -1 * image_in[554] -15 * image_in[555] -12 * image_in[556] +30 * image_in[557] +47 * image_in[558] +22 * image_in[559] +1 * image_in[560] -12 * image_in[561] +11 * image_in[562] +51 * image_in[563] +23 * image_in[564] -6 * image_in[565] +5 * image_in[566] +6 * image_in[567] -11 * image_in[568] +2 * image_in[569] -20 * image_in[570] +2 * image_in[571] -10 * image_in[572] -5 * image_in[573] +25 * image_in[574] +35 * image_in[575]
                            +44 * image_in[576] +46 * image_in[577] +37 * image_in[578] +38 * image_in[579] +39 * image_in[580] +7 * image_in[581] -9 * image_in[582] -4 * image_in[583] +42 * image_in[584] +33 * image_in[585] +33 * image_in[586] +6 * image_in[587] -2 * image_in[588] +10 * image_in[589] +45 * image_in[590] +59 * image_in[591] +23 * image_in[592] +14 * image_in[593] -6 * image_in[594] +2 * image_in[595] +5 * image_in[596] -5 * image_in[597] +5 * image_in[598] -16 * image_in[599] -7 * image_in[600] -2 * image_in[601] +10 * image_in[602] +15 * image_in[603] +36 * image_in[604] +34 * image_in[605] +41 * image_in[606] +45 * image_in[607]
                            +27 * image_in[608] +28 * image_in[609] +4 * image_in[610] +17 * image_in[611] +36 * image_in[612] +7 * image_in[613] +8 * image_in[614] -2 * image_in[615] +5 * image_in[616] -3 * image_in[617] +39 * image_in[618] +54 * image_in[619] +37 * image_in[620] +38 * image_in[621] +17 * image_in[622] -9 * image_in[623] +5 * image_in[624] +12 * image_in[625] +8 * image_in[626] -1 * image_in[627] -18 * image_in[628] -21 * image_in[629] -5 * image_in[630] +4 * image_in[631] +31 * image_in[633] +31 * image_in[634] +32 * image_in[635] +41 * image_in[636] +38 * image_in[637] +22 * image_in[638] +15 * image_in[639]
                            +21 * image_in[640] +7 * image_in[641] +17 * image_in[642] +6 * image_in[643] +20 * image_in[646] +36 * image_in[647] +25 * image_in[648] +28 * image_in[649] +22 * image_in[650] +14 * image_in[651] +7 * image_in[652] -1 * image_in[653] -9 * image_in[654] -2 * image_in[655] -10 * image_in[656] -12 * image_in[657] -18 * image_in[658] -7 * image_in[659] -13 * image_in[660] +18 * image_in[661] +40 * image_in[662] +33 * image_in[663] +47 * image_in[664] +33 * image_in[665] +37 * image_in[666] +22 * image_in[667] +15 * image_in[668] +1 * image_in[669] +23 * image_in[670] +2 * image_in[671]
                            +4 * image_in[672] +6 * image_in[673] +20 * image_in[674] +4 * image_in[675] +39 * image_in[676] +13 * image_in[677] +29 * image_in[678] +24 * image_in[679] +2 * image_in[680] +7 * image_in[681] +10 * image_in[682] -3 * image_in[683] -10 * image_in[684] -13 * image_in[685] -15 * image_in[686] -19 * image_in[687] -10 * image_in[688] +12 * image_in[689] +6 * image_in[690] +4 * image_in[691] +24 * image_in[692] +48 * image_in[693] +51 * image_in[694] +25 * image_in[695] +4 * image_in[696] +40 * image_in[697] +2 * image_in[698] -3 * image_in[699] +5 * image_in[700] -3 * image_in[701] -4 * image_in[702] -26 * image_in[703]
                            -11 * image_in[704] +27 * image_in[705] +25 * image_in[706] +12 * image_in[707] +25 * image_in[708] +21 * image_in[709] +21 * image_in[710] -2 * image_in[711] +11 * image_in[712] -1 * image_in[713] +3 * image_in[714] -38 * image_in[715] -24 * image_in[716] -30 * image_in[717] -16 * image_in[718] -10 * image_in[719] +22 * image_in[720] +5 * image_in[721] -11 * image_in[722] -8 * image_in[723] -22 * image_in[724] +2 * image_in[725] -1 * image_in[726] -3 * image_in[727] -3 * image_in[728] +6 * image_in[729] -4 * image_in[730] -1 * image_in[731] +29 * image_in[732] +28 * image_in[733] +36 * image_in[734] +24 * image_in[735]
                            +22 * image_in[736] +2 * image_in[737] +5 * image_in[738] -5 * image_in[739] -1 * image_in[740] -20 * image_in[741] +2 * image_in[742] -9 * image_in[743] +1 * image_in[744] -15 * image_in[745] +5 * image_in[746] -11 * image_in[747] +17 * image_in[748] +10 * image_in[749] -8 * image_in[750] +19 * image_in[751] -1 * image_in[752] -3 * image_in[753] +4 * image_in[754] +1 * image_in[755] +3 * image_in[757] -2 * image_in[758] +1 * image_in[759] +1 * image_in[760] -17 * image_in[761] -34 * image_in[762] -23 * image_in[763] -27 * image_in[764] -1 * image_in[765] -35 * image_in[766] -10 * image_in[767]
                            -8 * image_in[768] -35 * image_in[769] -14 * image_in[770] -1 * image_in[771] -4 * image_in[772] -35 * image_in[773] -33 * image_in[774] -11 * image_in[775] +2 * image_in[776] -6 * image_in[777] +16 * image_in[778] -4 * image_in[780] +1 * image_in[781] -2 * image_in[782];
                        if (layer1_out[4] < 0) layer1_out[4] = 0;
                        layer1_out[5] = -74 +5 * image_in[0] +5 * image_in[1] +2 * image_in[2] +1 * image_in[3] +5 * image_in[5] +4 * image_in[6] -4 * image_in[7] -6 * image_in[8] +2 * image_in[9] -4 * image_in[10] -2 * image_in[11] +6 * image_in[13] +6 * image_in[14] -5 * image_in[15] +4 * image_in[16] -2 * image_in[17] +3 * image_in[18] -6 * image_in[19] +5 * image_in[21] +5 * image_in[22] -3 * image_in[23] +6 * image_in[24] -4 * image_in[25] +4 * image_in[26] -4 * image_in[27] +4 * image_in[29] +6 * image_in[30] +4 * image_in[31]
                            +1 * image_in[32] -5 * image_in[33] +22 * image_in[34] +38 * image_in[35] +30 * image_in[36] +18 * image_in[37] +19 * image_in[38] +32 * image_in[39] +50 * image_in[40] +32 * image_in[41] -1 * image_in[42] +28 * image_in[43] +57 * image_in[44] +25 * image_in[45] +11 * image_in[46] +27 * image_in[47] +24 * image_in[48] +27 * image_in[49] +19 * image_in[50] +21 * image_in[51] +1 * image_in[52] -4 * image_in[53] -2 * image_in[54] -3 * image_in[55] -2 * image_in[56] +3 * image_in[57] +6 * image_in[58] -1 * image_in[59] +8 * image_in[60] +5 * image_in[61] +11 * image_in[62] +45 * image_in[63]
                            +44 * image_in[64] +61 * image_in[65] +66 * image_in[66] +59 * image_in[67] +58 * image_in[68] +33 * image_in[69] +28 * image_in[70] +16 * image_in[71] +37 * image_in[72] +18 * image_in[73] +22 * image_in[74] -4 * image_in[75] +22 * image_in[76] +31 * image_in[77] +16 * image_in[78] +34 * image_in[79] +36 * image_in[80] +25 * image_in[81] +3 * image_in[82] +4 * image_in[83] -3 * image_in[84] -6 * image_in[85] +17 * image_in[86] +4 * image_in[87] -5 * image_in[88] +21 * image_in[90] +30 * image_in[91] +56 * image_in[92] +81 * image_in[93] +68 * image_in[94] +97 * image_in[95]
                            +86 * image_in[96] +86 * image_in[97] +58 * image_in[98] +53 * image_in[99] +42 * image_in[100] +24 * image_in[101] +13 * image_in[102] -14 * image_in[103] -16 * image_in[104] -30 * image_in[105] -14 * image_in[106] +5 * image_in[107] +35 * image_in[108] -9 * image_in[109] +3 * image_in[110] -1 * image_in[111] +2 * image_in[112] -2 * image_in[113] -26 * image_in[114] +4 * image_in[115] -8 * image_in[116] +2 * image_in[117] +32 * image_in[118] +17 * image_in[119] +31 * image_in[120] +53 * image_in[121] +80 * image_in[122] +49 * image_in[123] +63 * image_in[124] +56 * image_in[125] +59 * image_in[126] +59 * image_in[127]
                            +39 * image_in[128] +50 * image_in[129] +41 * image_in[130] +6 * image_in[131] -6 * image_in[132] -58 * image_in[133] -45 * image_in[134] -47 * image_in[135] -76 * image_in[136] -7 * image_in[137] -9 * image_in[138] -5 * image_in[139] +2 * image_in[140] +2 * image_in[141] -3 * image_in[142] +19 * image_in[143] +12 * image_in[144] -32 * image_in[145] -12 * image_in[146] -5 * image_in[147] +4 * image_in[148] -1 * image_in[149] +19 * image_in[150] +17 * image_in[151] +31 * image_in[152] +47 * image_in[153] +39 * image_in[154] +37 * image_in[155] +31 * image_in[156] +30 * image_in[157] +37 * image_in[158] +12 * image_in[159]
                            +13 * image_in[160] +9 * image_in[161] -14 * image_in[162] -62 * image_in[163] -37 * image_in[164] -14 * image_in[165] +14 * image_in[166] -3 * image_in[167] +5 * image_in[168] -4 * image_in[169] -29 * image_in[170] +19 * image_in[171] -10 * image_in[172] -18 * image_in[173] -6 * image_in[174] +3 * image_in[175] -2 * image_in[176] +2 * image_in[178] +2 * image_in[179] +12 * image_in[180] +38 * image_in[181] +32 * image_in[182] +28 * image_in[183] +36 * image_in[184] +24 * image_in[185] +39 * image_in[186] +20 * image_in[187] +5 * image_in[188] +4 * image_in[189] -15 * image_in[190] -40 * image_in[191]
                            -71 * image_in[192] -28 * image_in[193] -38 * image_in[194] -4 * image_in[196] +32 * image_in[197] -7 * image_in[198] -7 * image_in[199] +28 * image_in[200] -8 * image_in[201] -2 * image_in[202] -17 * image_in[203] +2 * image_in[204] -7 * image_in[205] +7 * image_in[207] +20 * image_in[208] +20 * image_in[209] +32 * image_in[210] +32 * image_in[211] +31 * image_in[212] +16 * image_in[213] +24 * image_in[214] +10 * image_in[215] -7 * image_in[216] +1 * image_in[217] +1 * image_in[218] -32 * image_in[219] -33 * image_in[220] -52 * image_in[221] -30 * image_in[222] +5 * image_in[223]
                            -19 * image_in[224] -29 * image_in[225] -27 * image_in[226] +10 * image_in[227] +22 * image_in[228] -7 * image_in[229] +7 * image_in[230] -2 * image_in[231] -3 * image_in[232] +10 * image_in[233] +22 * image_in[234] +3 * image_in[235] +15 * image_in[236] +29 * image_in[237] +42 * image_in[238] +41 * image_in[239] +44 * image_in[240] +20 * image_in[241] +13 * image_in[242] +25 * image_in[243] +6 * image_in[244] +2 * image_in[245] +9 * image_in[246] -4 * image_in[247] -42 * image_in[248] -75 * image_in[249] -6 * image_in[250] +12 * image_in[251] -12 * image_in[252] -30 * image_in[253] -43 * image_in[254] +14 * image_in[255]
                            +30 * image_in[256] +12 * image_in[257] +13 * image_in[258] +14 * image_in[259] +15 * image_in[260] +13 * image_in[261] +17 * image_in[262] +11 * image_in[263] +2 * image_in[264] +28 * image_in[265] +52 * image_in[266] +28 * image_in[267] +20 * image_in[268] +16 * image_in[269] +24 * image_in[270] +13 * image_in[271] +1 * image_in[272] -12 * image_in[273] +9 * image_in[275] -17 * image_in[276] -65 * image_in[277] -21 * image_in[278] -18 * image_in[279] -20 * image_in[280] -33 * image_in[281] -12 * image_in[282] +8 * image_in[283] +25 * image_in[284] +20 * image_in[285] +34 * image_in[286] +10 * image_in[287]
                            +2 * image_in[288] +9 * image_in[289] +5 * image_in[290] +4 * image_in[291] +6 * image_in[292] +16 * image_in[293] +38 * image_in[294] -5 * image_in[295] +2 * image_in[296] +17 * image_in[297] +27 * image_in[298] +5 * image_in[299] +17 * image_in[300] +8 * image_in[301] +29 * image_in[302] +61 * image_in[303] +37 * image_in[304] -71 * image_in[305] -8 * image_in[306] +10 * image_in[307] -19 * image_in[308] -21 * image_in[309] -23 * image_in[310] +24 * image_in[312] +14 * image_in[313] -5 * image_in[314] +2 * image_in[315] +6 * image_in[316] -21 * image_in[317] -26 * image_in[318] -7 * image_in[319]
                            -40 * image_in[320] +11 * image_in[321] +9 * image_in[322] -38 * image_in[323] -41 * image_in[324] -23 * image_in[325] -1 * image_in[326] +24 * image_in[327] +31 * image_in[328] +27 * image_in[329] +38 * image_in[330] +73 * image_in[331] +57 * image_in[332] +1 * image_in[333] -32 * image_in[334] -19 * image_in[335] -18 * image_in[336] -31 * image_in[337] -23 * image_in[338] -5 * image_in[339] +4 * image_in[340] +2 * image_in[341] -12 * image_in[342] -19 * image_in[343] -30 * image_in[344] -14 * image_in[345] -24 * image_in[346] -35 * image_in[347] -16 * image_in[348] +10 * image_in[349] -8 * image_in[350] -31 * image_in[351]
                            -45 * image_in[352] -12 * image_in[353] +2 * image_in[354] +20 * image_in[355] +24 * image_in[356] +18 * image_in[357] +45 * image_in[358] +75 * image_in[359] +94 * image_in[360] +42 * image_in[361] +24 * image_in[362] -21 * image_in[363] -4 * image_in[364] -12 * image_in[365] -18 * image_in[366] +18 * image_in[367] -55 * image_in[368] -34 * image_in[369] -27 * image_in[370] -32 * image_in[371] -9 * image_in[372] -8 * image_in[373] -14 * image_in[374] -3 * image_in[375] +10 * image_in[376] +28 * image_in[377] -4 * image_in[378] -28 * image_in[379] -24 * image_in[380] -18 * image_in[381] -17 * image_in[382] +11 * image_in[383]
                            -6 * image_in[384] +17 * image_in[385] +36 * image_in[386] +68 * image_in[387] +73 * image_in[388] +59 * image_in[389] +22 * image_in[390] +34 * image_in[391] +6 * image_in[392] -6 * image_in[393] -27 * image_in[394] +2 * image_in[395] -58 * image_in[396] -25 * image_in[397] -10 * image_in[398] -1 * image_in[399] -2 * image_in[400] -4 * image_in[401] +7 * image_in[403] +24 * image_in[404] +24 * image_in[405] -8 * image_in[406] -10 * image_in[407] -39 * image_in[408] -30 * image_in[409] -17 * image_in[410] -18 * image_in[411] -3 * image_in[412] +19 * image_in[413] +9 * image_in[414] +35 * image_in[415]
                            +54 * image_in[416] +41 * image_in[417] +53 * image_in[418] -5 * image_in[419] -3 * image_in[420] -13 * image_in[421] -46 * image_in[422] -17 * image_in[423] +3 * image_in[424] +14 * image_in[425] +2 * image_in[426] +14 * image_in[427] +7 * image_in[428] +9 * image_in[429] +21 * image_in[430] +16 * image_in[431] +18 * image_in[432] +22 * image_in[433] -8 * image_in[434] -32 * image_in[435] -30 * image_in[436] -28 * image_in[437] -15 * image_in[438] +9 * image_in[440] +5 * image_in[441] +1 * image_in[442] +20 * image_in[443] +68 * image_in[444] +64 * image_in[445] +39 * image_in[446] +13 * image_in[447]
                            +1 * image_in[448] -5 * image_in[449] +3 * image_in[450] +22 * image_in[451] +21 * image_in[452] +24 * image_in[453] +11 * image_in[454] +14 * image_in[455] +4 * image_in[456] +32 * image_in[457] +43 * image_in[458] +42 * image_in[459] +24 * image_in[460] -8 * image_in[461] -10 * image_in[462] -39 * image_in[463] -31 * image_in[464] -8 * image_in[465] -7 * image_in[466] -6 * image_in[467] +1 * image_in[468] +24 * image_in[469] +13 * image_in[470] +31 * image_in[471] +37 * image_in[472] +63 * image_in[473] +44 * image_in[474] +29 * image_in[475] -5 * image_in[476] -12 * image_in[477] +34 * image_in[479]
                            +15 * image_in[480] +23 * image_in[481] +24 * image_in[482] +19 * image_in[483] +22 * image_in[484] +37 * image_in[485] +61 * image_in[486] +46 * image_in[487] +20 * image_in[488] -16 * image_in[489] -43 * image_in[490] -28 * image_in[491] -17 * image_in[492] -10 * image_in[493] -5 * image_in[494] +18 * image_in[495] -4 * image_in[496] -9 * image_in[497] +29 * image_in[498] +30 * image_in[499] +34 * image_in[500] +71 * image_in[501] +53 * image_in[502] -1 * image_in[503] -2 * image_in[504] -8 * image_in[505] +14 * image_in[506] +7 * image_in[507] +6 * image_in[508] +18 * image_in[509] +17 * image_in[510] +29 * image_in[511]
                            +35 * image_in[512] +49 * image_in[513] +69 * image_in[514] +37 * image_in[515] +21 * image_in[516] -15 * image_in[517] -29 * image_in[518] -6 * image_in[519] +11 * image_in[520] +25 * image_in[521] +22 * image_in[522] +31 * image_in[523] +7 * image_in[524] +11 * image_in[525] +36 * image_in[526] +47 * image_in[527] +69 * image_in[528] +75 * image_in[529] +32 * image_in[530] +37 * image_in[531] +5 * image_in[532] -5 * image_in[533] -14 * image_in[534] -8 * image_in[535] +10 * image_in[536] +10 * image_in[537] +22 * image_in[538] +42 * image_in[539] +37 * image_in[540] +53 * image_in[541] +70 * image_in[542] +44 * image_in[543]
                            +40 * image_in[544] +24 * image_in[545] +7 * image_in[546] +15 * image_in[547] +15 * image_in[548] +36 * image_in[549] +33 * image_in[550] +27 * image_in[551] +45 * image_in[552] +40 * image_in[553] +62 * image_in[554] +48 * image_in[555] +17 * image_in[556] +53 * image_in[557] +42 * image_in[558] +15 * image_in[559] +2 * image_in[560] +17 * image_in[561] -13 * image_in[562] +2 * image_in[563] +34 * image_in[564] +40 * image_in[565] +38 * image_in[566] +57 * image_in[567] +60 * image_in[568] +43 * image_in[569] +63 * image_in[570] +41 * image_in[571] +54 * image_in[572] +42 * image_in[573] +23 * image_in[574] +19 * image_in[575]
                            +19 * image_in[576] +15 * image_in[577] +36 * image_in[578] +32 * image_in[579] +40 * image_in[580] +59 * image_in[581] +23 * image_in[582] +27 * image_in[583] +27 * image_in[585] +8 * image_in[586] +4 * image_in[588] +14 * image_in[589] +23 * image_in[590] +46 * image_in[591] +29 * image_in[592] +27 * image_in[593] +33 * image_in[594] +46 * image_in[595] +26 * image_in[596] +30 * image_in[597] +29 * image_in[598] +55 * image_in[599] +41 * image_in[600] +49 * image_in[601] +50 * image_in[602] +34 * image_in[603] +30 * image_in[604] +24 * image_in[605] +42 * image_in[606] +37 * image_in[607]
                            +21 * image_in[608] +21 * image_in[609] +28 * image_in[610] +38 * image_in[611] +7 * image_in[612] +34 * image_in[613] +8 * image_in[614] -4 * image_in[615] -5 * image_in[616] +6 * image_in[617] +38 * image_in[618] +58 * image_in[619] -1 * image_in[620] +1 * image_in[621] +46 * image_in[622] +26 * image_in[623] +36 * image_in[624] +41 * image_in[625] +34 * image_in[626] +39 * image_in[627] +41 * image_in[628] +45 * image_in[629] +29 * image_in[630] +35 * image_in[631] +30 * image_in[632] +15 * image_in[633] +29 * image_in[634] +16 * image_in[635] +25 * image_in[636] -3 * image_in[637] +15 * image_in[638] -1 * image_in[639] +10 * image_in[641] -5 * image_in[642] -3 * image_in[643] -6 * image_in[644] +2 * image_in[645] +22 * image_in[646] +27 * image_in[647] -20 * image_in[648] -12 * image_in[649] -12 * image_in[650] -3 * image_in[651] +35 * image_in[652] +20 * image_in[653] +29 * image_in[654] +26 * image_in[655] +41 * image_in[656] +33 * image_in[657] +24 * image_in[658] +13 * image_in[659] -2 * image_in[660] -1 * image_in[661] +5 * image_in[662] +9 * image_in[663] +8 * image_in[664] -1 * image_in[665] +21 * image_in[666] +25 * image_in[667] +17 * image_in[668] +1 * image_in[669] -20 * image_in[670] -1 * image_in[671]
                            -6 * image_in[672] -1 * image_in[673] +17 * image_in[674] -33 * image_in[675] -5 * image_in[676] -52 * image_in[677] -35 * image_in[678] -39 * image_in[679] -36 * image_in[680] -2 * image_in[681] -11 * image_in[682] -10 * image_in[683] +14 * image_in[684] -1 * image_in[685] +13 * image_in[686] +9 * image_in[687] +12 * image_in[688] +14 * image_in[689] +18 * image_in[690] +1 * image_in[691] -14 * image_in[692] +13 * image_in[693] -19 * image_in[694] -17 * image_in[695] +23 * image_in[696] +39 * image_in[697] +5 * image_in[698] -2 * image_in[699] +6 * image_in[700] -2 * image_in[701] -24 * image_in[703]
                            -30 * image_in[704] -26 * image_in[705] -1 * image_in[706] -19 * image_in[707] -11 * image_in[708] -31 * image_in[709] -25 * image_in[710] -21 * image_in[711] -8 * image_in[713] -6 * image_in[714] +11 * image_in[715] +26 * image_in[716] +19 * image_in[717] +11 * image_in[718] +16 * image_in[719] +14 * image_in[720] +5 * image_in[721] -7 * image_in[722] -17 * image_in[723] +4 * image_in[724] +2 * image_in[726] -2 * image_in[727] -2 * image_in[728] -6 * image_in[729] +4 * image_in[730] +15 * image_in[732] -6 * image_in[733] +4 * image_in[734] +5 * image_in[735]
                            +7 * image_in[736] -1 * image_in[737] +9 * image_in[738] +14 * image_in[739] +29 * image_in[740] +2 * image_in[741] +9 * image_in[742] +6 * image_in[743] +17 * image_in[744] +18 * image_in[745] +25 * image_in[746] +24 * image_in[747] +17 * image_in[748] +21 * image_in[749] +7 * image_in[750] +21 * image_in[751] -6 * image_in[752] -4 * image_in[753] -4 * image_in[754] +4 * image_in[755] +2 * image_in[756] -5 * image_in[757] +5 * image_in[758] +5 * image_in[759] -4 * image_in[760] -20 * image_in[761] -34 * image_in[762] -51 * image_in[763] -15 * image_in[764] +4 * image_in[765] -3 * image_in[766] +24 * image_in[767]
                            +17 * image_in[768] -25 * image_in[769] +14 * image_in[770] -9 * image_in[771] -17 * image_in[772] -36 * image_in[773] -43 * image_in[774] +11 * image_in[775] -4 * image_in[776] +14 * image_in[777] -19 * image_in[778] +2 * image_in[779] +4 * image_in[780] +5 * image_in[781] +5 * image_in[782] -1 * image_in[783];
                        if (layer1_out[5] < 0) layer1_out[5] = 0;
                        layer1_out[6] = 70 +5 * image_in[0] +2 * image_in[3] +3 * image_in[4] -4 * image_in[5] -4 * image_in[6] -1 * image_in[7] +5 * image_in[8] -6 * image_in[9] -3 * image_in[10] +4 * image_in[11] +2 * image_in[12] -8 * image_in[13] -8 * image_in[14] +4 * image_in[15] +3 * image_in[16] -4 * image_in[17] -1 * image_in[18] -4 * image_in[19] +3 * image_in[20] +6 * image_in[21] -6 * image_in[22] +2 * image_in[24] -5 * image_in[25] -6 * image_in[26] -2 * image_in[27] -1 * image_in[28] -1 * image_in[29] +5 * image_in[31]
                            +5 * image_in[32] +6 * image_in[33] -22 * image_in[34] -31 * image_in[35] -22 * image_in[36] -14 * image_in[37] -22 * image_in[38] -2 * image_in[39] -20 * image_in[40] -45 * image_in[41] -8 * image_in[42] -47 * image_in[43] -35 * image_in[44] -38 * image_in[45] -31 * image_in[46] -32 * image_in[47] -30 * image_in[48] -16 * image_in[49] -27 * image_in[50] -14 * image_in[51] -3 * image_in[52] +2 * image_in[53] +5 * image_in[55] -4 * image_in[56] +5 * image_in[57] +1 * image_in[58] +6 * image_in[59] -6 * image_in[60] +5 * image_in[61] -33 * image_in[62] -40 * image_in[63]
                            -50 * image_in[64] -66 * image_in[65] -73 * image_in[66] -62 * image_in[67] -42 * image_in[68] -48 * image_in[69] -65 * image_in[70] -66 * image_in[71] -61 * image_in[72] -28 * image_in[73] -5 * image_in[74] -10 * image_in[75] -48 * image_in[76] -35 * image_in[77] -39 * image_in[78] -33 * image_in[79] -39 * image_in[80] -18 * image_in[81] +2 * image_in[82] +6 * image_in[83] +1 * image_in[84] +3 * image_in[85] -17 * image_in[86] +2 * image_in[87] -1 * image_in[88] +24 * image_in[89] -26 * image_in[90] -16 * image_in[91] +5 * image_in[92] -36 * image_in[93] -23 * image_in[94] -5 * image_in[95]
                            -10 * image_in[96] -24 * image_in[97] +5 * image_in[98] -13 * image_in[99] -18 * image_in[100] +1 * image_in[101] +13 * image_in[102] +19 * image_in[103] +28 * image_in[104] +6 * image_in[105] +1 * image_in[106] -8 * image_in[107] -15 * image_in[108] +23 * image_in[109] -2 * image_in[110] +1 * image_in[111] +3 * image_in[112] +2 * image_in[113] -16 * image_in[114] -4 * image_in[115] +10 * image_in[116] -1 * image_in[117] -25 * image_in[118] -6 * image_in[120] -15 * image_in[121] -15 * image_in[122] +4 * image_in[123] -6 * image_in[124] -25 * image_in[125] -13 * image_in[126] +2 * image_in[127]
                            +6 * image_in[128] +7 * image_in[129] +12 * image_in[130] +9 * image_in[131] -1 * image_in[132] +34 * image_in[133] +19 * image_in[134] +23 * image_in[135] +65 * image_in[136] +31 * image_in[137] +20 * image_in[138] -4 * image_in[139] -1 * image_in[140] +3 * image_in[141] +3 * image_in[142] -14 * image_in[144] +6 * image_in[145] +14 * image_in[146] +14 * image_in[147] +6 * image_in[148] +16 * image_in[149] -5 * image_in[150] +4 * image_in[151] -23 * image_in[152] -19 * image_in[153] -16 * image_in[154] -2 * image_in[155] +6 * image_in[156] +14 * image_in[157] +11 * image_in[158] +7 * image_in[159]
                            +11 * image_in[160] -13 * image_in[161] +3 * image_in[162] +18 * image_in[163] +7 * image_in[164] +42 * image_in[165] +2 * image_in[166] +3 * image_in[167] +1 * image_in[168] -3 * image_in[169] +16 * image_in[170] +35 * image_in[172] +5 * image_in[173] +23 * image_in[174] +3 * image_in[175] +20 * image_in[176] +11 * image_in[177] +12 * image_in[178] -3 * image_in[179] +5 * image_in[180] -7 * image_in[181] +7 * image_in[182] +8 * image_in[183] +12 * image_in[184] +16 * image_in[185] +16 * image_in[186] +17 * image_in[187] +8 * image_in[188] +17 * image_in[189] +14 * image_in[190] +15 * image_in[191]
                            +49 * image_in[192] +42 * image_in[193] +34 * image_in[194] -12 * image_in[195] -2 * image_in[196] +37 * image_in[197] -8 * image_in[198] +19 * image_in[199] -7 * image_in[200] +21 * image_in[201] +13 * image_in[202] +25 * image_in[203] +15 * image_in[204] +27 * image_in[205] +10 * image_in[206] +2 * image_in[207] +7 * image_in[208] +12 * image_in[209] +15 * image_in[210] +20 * image_in[211] +13 * image_in[212] +44 * image_in[213] +23 * image_in[214] +30 * image_in[215] +15 * image_in[216] +13 * image_in[217] +7 * image_in[218] +37 * image_in[219] +59 * image_in[220] +70 * image_in[221] +27 * image_in[222] -2 * image_in[223]
                            +2 * image_in[224] +13 * image_in[225] +23 * image_in[226] +1 * image_in[227] -9 * image_in[228] +15 * image_in[229] +14 * image_in[230] -3 * image_in[231] +4 * image_in[232] +24 * image_in[233] +15 * image_in[234] +18 * image_in[235] -3 * image_in[236] +9 * image_in[237] +4 * image_in[238] +12 * image_in[239] +28 * image_in[240] +38 * image_in[241] +49 * image_in[242] +32 * image_in[243] +41 * image_in[244] +32 * image_in[245] +38 * image_in[246] +51 * image_in[247] +93 * image_in[248] +88 * image_in[249] +40 * image_in[250] +5 * image_in[251] +2 * image_in[252] +14 * image_in[253] +28 * image_in[254] +7 * image_in[255]
                            -8 * image_in[256] +4 * image_in[257] -10 * image_in[258] +6 * image_in[259] +10 * image_in[260] +15 * image_in[261] +8 * image_in[262] +4 * image_in[263] +8 * image_in[264] +16 * image_in[265] +6 * image_in[266] -1 * image_in[267] +17 * image_in[268] +35 * image_in[269] +47 * image_in[270] +38 * image_in[271] +38 * image_in[272] +50 * image_in[273] +57 * image_in[274] +63 * image_in[275] +98 * image_in[276] +100 * image_in[277] +36 * image_in[278] +15 * image_in[279] +10 * image_in[280] -16 * image_in[281] +21 * image_in[282] +24 * image_in[283] -6 * image_in[284] -12 * image_in[285] -11 * image_in[286] +14 * image_in[287]
                            -4 * image_in[288] +15 * image_in[289] -4 * image_in[290] -3 * image_in[291] +9 * image_in[292] +11 * image_in[293] +6 * image_in[294] +14 * image_in[295] +30 * image_in[296] +32 * image_in[297] +28 * image_in[298] +19 * image_in[299] +40 * image_in[300] +37 * image_in[301] +37 * image_in[302] +61 * image_in[303] +106 * image_in[304] +127 * image_in[305] +64 * image_in[306] +18 * image_in[307] +7 * image_in[308] -3 * image_in[309] +17 * image_in[310] +28 * image_in[311] -13 * image_in[312] -28 * image_in[313] +12 * image_in[314] -10 * image_in[315] +4 * image_in[316] +12 * image_in[317] +14 * image_in[318] +24 * image_in[319]
                            +35 * image_in[320] +23 * image_in[321] +10 * image_in[322] +13 * image_in[323] +5 * image_in[324] +32 * image_in[325] +19 * image_in[326] +11 * image_in[327] -12 * image_in[328] -15 * image_in[329] -5 * image_in[330] -1 * image_in[331] +41 * image_in[332] +74 * image_in[333] +53 * image_in[334] -16 * image_in[335] +4 * image_in[336] -4 * image_in[337] +12 * image_in[338] +15 * image_in[339] -16 * image_in[340] -25 * image_in[341] +13 * image_in[342] +12 * image_in[344] +17 * image_in[345] +45 * image_in[346] +41 * image_in[347] +41 * image_in[348] +23 * image_in[349] -6 * image_in[350] +2 * image_in[351] +13 * image_in[353] +4 * image_in[354] -6 * image_in[355] -27 * image_in[356] -31 * image_in[357] -52 * image_in[358] -72 * image_in[359] -58 * image_in[360] +13 * image_in[361] +1 * image_in[362] -19 * image_in[363] +4 * image_in[364] -1 * image_in[365] -5 * image_in[366] +16 * image_in[368] +24 * image_in[369] +22 * image_in[370] +31 * image_in[371] +17 * image_in[372] +26 * image_in[373] +54 * image_in[374] +57 * image_in[375] +26 * image_in[376] +19 * image_in[377] -9 * image_in[378] -17 * image_in[379] -2 * image_in[380] +12 * image_in[381] +27 * image_in[382] +6 * image_in[383]
                            -1 * image_in[384] -16 * image_in[385] -14 * image_in[386] -59 * image_in[387] -52 * image_in[388] -34 * image_in[389] -24 * image_in[390] -31 * image_in[391] -2 * image_in[392] -23 * image_in[393] -2 * image_in[395] +51 * image_in[396] +14 * image_in[397] +4 * image_in[399] +10 * image_in[400] +31 * image_in[401] +47 * image_in[402] +26 * image_in[403] +11 * image_in[404] -12 * image_in[405] -14 * image_in[406] -19 * image_in[407] -10 * image_in[408] +40 * image_in[409] +33 * image_in[410] +22 * image_in[411] +9 * image_in[412] +14 * image_in[413] +16 * image_in[414] -1 * image_in[415]
                            -13 * image_in[416] -55 * image_in[417] -55 * image_in[418] -3 * image_in[419] +4 * image_in[420] +22 * image_in[421] +34 * image_in[422] -11 * image_in[423] +19 * image_in[424] +7 * image_in[425] -1 * image_in[426] -5 * image_in[427] -1 * image_in[428] +13 * image_in[429] +26 * image_in[430] +14 * image_in[431] +1 * image_in[432] -26 * image_in[433] -38 * image_in[434] -8 * image_in[435] +4 * image_in[436] +36 * image_in[437] +37 * image_in[438] +31 * image_in[439] +31 * image_in[440] +28 * image_in[441] +34 * image_in[442] +50 * image_in[443] -21 * image_in[444] -75 * image_in[445] -34 * image_in[446] -23 * image_in[447]
                            +1 * image_in[448] +3 * image_in[449] +27 * image_in[450] -29 * image_in[451] -8 * image_in[452] +4 * image_in[453] -3 * image_in[454] -6 * image_in[455] -4 * image_in[456] -23 * image_in[457] -21 * image_in[458] -22 * image_in[459] -9 * image_in[460] -15 * image_in[461] -28 * image_in[462] -4 * image_in[463] +10 * image_in[464] +40 * image_in[465] +43 * image_in[466] +42 * image_in[467] +39 * image_in[468] +20 * image_in[469] +38 * image_in[470] +30 * image_in[471] -3 * image_in[472] -89 * image_in[473] -62 * image_in[474] -34 * image_in[475] -3 * image_in[476] +5 * image_in[477] -10 * image_in[478] -7 * image_in[479]
                            +14 * image_in[480] +24 * image_in[481] +32 * image_in[482] +5 * image_in[483] -10 * image_in[484] -35 * image_in[485] -42 * image_in[486] -44 * image_in[487] -41 * image_in[488] -35 * image_in[489] -14 * image_in[490] +12 * image_in[491] +29 * image_in[492] +48 * image_in[493] +44 * image_in[494] +34 * image_in[495] +23 * image_in[496] +22 * image_in[497] +8 * image_in[498] +6 * image_in[499] -18 * image_in[500] -90 * image_in[501] -56 * image_in[502] -1 * image_in[503] -6 * image_in[504] +7 * image_in[505] -3 * image_in[506] +22 * image_in[507] +23 * image_in[508] +38 * image_in[509] +54 * image_in[510] +19 * image_in[511] -29 * image_in[513] -28 * image_in[514] -27 * image_in[515] -21 * image_in[516] -14 * image_in[517] -9 * image_in[518] +21 * image_in[519] +27 * image_in[520] +30 * image_in[521] +8 * image_in[522] +11 * image_in[523] +10 * image_in[524] +14 * image_in[525] +8 * image_in[526] -31 * image_in[527] -54 * image_in[528] -86 * image_in[529] -37 * image_in[530] -18 * image_in[531] -1 * image_in[532] +5 * image_in[533] +20 * image_in[534] +47 * image_in[535] +14 * image_in[536] +54 * image_in[537] +28 * image_in[538] +13 * image_in[539] +16 * image_in[540] -3 * image_in[541] -15 * image_in[542] -15 * image_in[543]
                            -2 * image_in[544] -10 * image_in[545] +3 * image_in[546] +13 * image_in[547] +4 * image_in[548] +12 * image_in[549] +2 * image_in[550] -9 * image_in[551] -12 * image_in[552] -3 * image_in[553] -28 * image_in[554] -24 * image_in[555] -13 * image_in[556] -42 * image_in[557] -44 * image_in[558] -11 * image_in[559] +3 * image_in[560] +23 * image_in[561] +16 * image_in[562] +17 * image_in[563] +12 * image_in[564] +27 * image_in[565] +18 * image_in[566] -5 * image_in[567] +3 * image_in[568] +6 * image_in[569] -7 * image_in[570] -8 * image_in[572] +6 * image_in[573] +9 * image_in[574] +6 * image_in[575]
                            -2 * image_in[576] -2 * image_in[577] -15 * image_in[578] -16 * image_in[579] -22 * image_in[580] -28 * image_in[581] -8 * image_in[582] -18 * image_in[583] -39 * image_in[584] -25 * image_in[585] -23 * image_in[586] -2 * image_in[587] +7 * image_in[589] -4 * image_in[590] -6 * image_in[591] -8 * image_in[592] -7 * image_in[593] -2 * image_in[594] -8 * image_in[595] +5 * image_in[596] +4 * image_in[597] -3 * image_in[598] +1 * image_in[599] +11 * image_in[600] +1 * image_in[601] +2 * image_in[602] -2 * image_in[604] -22 * image_in[605] -29 * image_in[606] -41 * image_in[607]
                            -28 * image_in[608] -25 * image_in[609] -14 * image_in[610] -32 * image_in[611] -40 * image_in[612] -22 * image_in[613] -2 * image_in[614] +5 * image_in[615] +3 * image_in[616] -6 * image_in[617] +8 * image_in[618] +3 * image_in[619] -7 * image_in[620] -45 * image_in[621] -31 * image_in[622] +5 * image_in[623] +5 * image_in[624] +6 * image_in[625] +4 * image_in[626] +16 * image_in[627] +19 * image_in[628] +30 * image_in[629] +3 * image_in[630] +5 * image_in[631] +8 * image_in[632] -15 * image_in[633] -28 * image_in[634] -24 * image_in[635] -32 * image_in[636] -22 * image_in[637] -14 * image_in[638] -4 * image_in[639]
                            -19 * image_in[640] -11 * image_in[641] -12 * image_in[642] +3 * image_in[645] +17 * image_in[646] +46 * image_in[647] +24 * image_in[648] +2 * image_in[649] +11 * image_in[650] +18 * image_in[651] +9 * image_in[652] +26 * image_in[653] +41 * image_in[654] +31 * image_in[655] +14 * image_in[656] +11 * image_in[657] +28 * image_in[658] +1 * image_in[659] -12 * image_in[661] -16 * image_in[662] -22 * image_in[663] -18 * image_in[664] -20 * image_in[665] -35 * image_in[666] -12 * image_in[667] +4 * image_in[668] +4 * image_in[669] -16 * image_in[670] -2 * image_in[671]
                            -1 * image_in[672] +6 * image_in[673] +18 * image_in[674] +54 * image_in[675] +62 * image_in[676] +41 * image_in[677] +38 * image_in[678] +63 * image_in[679] +34 * image_in[680] +29 * image_in[681] +39 * image_in[682] +47 * image_in[683] +30 * image_in[684] +46 * image_in[685] +35 * image_in[686] +29 * image_in[687] +23 * image_in[688] +12 * image_in[689] -26 * image_in[690] -30 * image_in[691] -14 * image_in[692] -26 * image_in[693] +11 * image_in[694] +22 * image_in[695] -33 * image_in[697] -3 * image_in[698] +5 * image_in[699] +4 * image_in[700] -6 * image_in[701] -4 * image_in[702] +33 * image_in[703]
                            +65 * image_in[704] +81 * image_in[705] +73 * image_in[706] +69 * image_in[707] +69 * image_in[708] +80 * image_in[709] +88 * image_in[710] +79 * image_in[711] +69 * image_in[712] +74 * image_in[713] +35 * image_in[714] +51 * image_in[715] +36 * image_in[716] +28 * image_in[717] +20 * image_in[718] +23 * image_in[719] -11 * image_in[720] +11 * image_in[721] +50 * image_in[722] +40 * image_in[723] +26 * image_in[724] -5 * image_in[725] -1 * image_in[726] +3 * image_in[727] -4 * image_in[728] +2 * image_in[729] +4 * image_in[730] +4 * image_in[731] -22 * image_in[732] -19 * image_in[733] -2 * image_in[734] -7 * image_in[735]
                            -13 * image_in[736] +11 * image_in[737] +18 * image_in[738] +24 * image_in[739] +26 * image_in[740] +40 * image_in[741] +9 * image_in[742] +26 * image_in[743] +38 * image_in[744] +11 * image_in[745] +9 * image_in[746] +13 * image_in[748] +7 * image_in[749] -3 * image_in[750] -18 * image_in[751] -6 * image_in[752] +1 * image_in[753] -2 * image_in[754] +1 * image_in[755] -3 * image_in[756] +4 * image_in[757] -3 * image_in[758] -5 * image_in[759] +4 * image_in[760] +22 * image_in[761] +30 * image_in[762] -20 * image_in[763] -10 * image_in[764] -5 * image_in[765] +10 * image_in[766]
                            +4 * image_in[768] +15 * image_in[769] -22 * image_in[770] -17 * image_in[771] -15 * image_in[772] +11 * image_in[773] +23 * image_in[774] -12 * image_in[775] -5 * image_in[776] -13 * image_in[777] -7 * image_in[778] -1 * image_in[780] -1 * image_in[781] -5 * image_in[782];
                        if (layer1_out[6] < 0) layer1_out[6] = 0;
                        layer1_out[7] = 127 +6 * image_in[0] +1 * image_in[1] +1 * image_in[2] +1 * image_in[3] +3 * image_in[4] -6 * image_in[5] +2 * image_in[6] +1 * image_in[7] -4 * image_in[8] -2 * image_in[9] -4 * image_in[10] -5 * image_in[11] +11 * image_in[13] -4 * image_in[14] -2 * image_in[15] -4 * image_in[16] -5 * image_in[17] -2 * image_in[18] -4 * image_in[19] +2 * image_in[20] +2 * image_in[21] -4 * image_in[22] +4 * image_in[24] +3 * image_in[25] -3 * image_in[26] -3 * image_in[27] -4 * image_in[28] -2 * image_in[29] -5 * image_in[30] -5 * image_in[31]
                            +5 * image_in[32] -3 * image_in[33] +7 * image_in[34] +27 * image_in[35] +22 * image_in[36] +22 * image_in[37] +19 * image_in[38] +38 * image_in[39] +48 * image_in[40] +51 * image_in[41] +13 * image_in[42] +15 * image_in[43] +13 * image_in[44] +21 * image_in[45] +27 * image_in[46] +21 * image_in[47] +27 * image_in[48] +13 * image_in[49] +11 * image_in[50] +12 * image_in[51] +4 * image_in[52] -6 * image_in[53] -4 * image_in[54] +2 * image_in[55] +3 * image_in[56] -4 * image_in[58] -6 * image_in[59] +8 * image_in[60] +3 * image_in[61] +22 * image_in[62] +38 * image_in[63]
                            +34 * image_in[64] +13 * image_in[65] +44 * image_in[66] +15 * image_in[67] +21 * image_in[68] -5 * image_in[69] +5 * image_in[70] +7 * image_in[71] -1 * image_in[72] +10 * image_in[73] +23 * image_in[74] +29 * image_in[75] +38 * image_in[76] +28 * image_in[77] +32 * image_in[78] +31 * image_in[79] -5 * image_in[80] -12 * image_in[81] +1 * image_in[82] -1 * image_in[83] +2 * image_in[84] -3 * image_in[85] +7 * image_in[86] -5 * image_in[87] +5 * image_in[88] -26 * image_in[89] -3 * image_in[90] -5 * image_in[91] -5 * image_in[92] +12 * image_in[93] -8 * image_in[94] -7 * image_in[95]
                            -7 * image_in[96] +16 * image_in[97] -6 * image_in[98] +7 * image_in[99] +4 * image_in[100] +7 * image_in[101] +11 * image_in[102] +24 * image_in[103] +26 * image_in[104] +47 * image_in[105] +46 * image_in[106] +31 * image_in[107] +36 * image_in[108] +3 * image_in[110] +1 * image_in[111] +1 * image_in[112] -5 * image_in[113] -4 * image_in[114] -1 * image_in[115] +6 * image_in[116] -33 * image_in[117] -44 * image_in[118] -20 * image_in[119] -27 * image_in[120] -21 * image_in[121] -22 * image_in[122] -6 * image_in[123] -19 * image_in[124] -16 * image_in[125] -6 * image_in[126] +1 * image_in[127]
                            -1 * image_in[128] +24 * image_in[129] +7 * image_in[130] +14 * image_in[131] +5 * image_in[132] +36 * image_in[133] +39 * image_in[134] +65 * image_in[135] +35 * image_in[136] +18 * image_in[137] -9 * image_in[138] -6 * image_in[139] -2 * image_in[140] -3 * image_in[141] -1 * image_in[142] -21 * image_in[143] -44 * image_in[144] -63 * image_in[145] -26 * image_in[146] -32 * image_in[147] -4 * image_in[148] -3 * image_in[149] +24 * image_in[150] +14 * image_in[151] -7 * image_in[152] -2 * image_in[153] +2 * image_in[154] -7 * image_in[155] -5 * image_in[156] +17 * image_in[157] +38 * image_in[158] +6 * image_in[159]
                            +25 * image_in[160] +20 * image_in[161] +24 * image_in[162] +34 * image_in[163] +45 * image_in[164] +20 * image_in[165] +8 * image_in[166] -4 * image_in[167] -5 * image_in[168] -4 * image_in[169] -3 * image_in[170] -36 * image_in[171] -26 * image_in[172] -20 * image_in[173] -30 * image_in[174] +8 * image_in[175] -5 * image_in[176] +2 * image_in[177] +3 * image_in[178] +19 * image_in[179] +25 * image_in[180] +2 * image_in[181] +10 * image_in[182] -5 * image_in[183] -3 * image_in[184] +10 * image_in[185] +18 * image_in[186] +15 * image_in[187] +12 * image_in[188] +21 * image_in[189] +23 * image_in[190] +19 * image_in[191]
                            +49 * image_in[192] +15 * image_in[193] +20 * image_in[194] +5 * image_in[195] -2 * image_in[196] -25 * image_in[197] +9 * image_in[198] -31 * image_in[199] -50 * image_in[200] -28 * image_in[201] -12 * image_in[202] +15 * image_in[203] +20 * image_in[204] +31 * image_in[205] +28 * image_in[206] +50 * image_in[207] +35 * image_in[208] +25 * image_in[209] +14 * image_in[210] +4 * image_in[211] +4 * image_in[212] +19 * image_in[213] +25 * image_in[214] +22 * image_in[215] +20 * image_in[216] +16 * image_in[217] +32 * image_in[218] +32 * image_in[219] +49 * image_in[220] +39 * image_in[221] +29 * image_in[222] -10 * image_in[223]
                            -3 * image_in[224] -2 * image_in[225] +5 * image_in[226] -33 * image_in[227] -64 * image_in[228] -29 * image_in[229] -17 * image_in[230] -4 * image_in[231] +14 * image_in[232] +23 * image_in[233] +24 * image_in[234] +41 * image_in[235] +22 * image_in[236] +13 * image_in[237] -8 * image_in[238] -8 * image_in[239] +6 * image_in[240] +19 * image_in[241] +7 * image_in[242] +19 * image_in[243] +21 * image_in[244] +13 * image_in[245] +5 * image_in[246] +38 * image_in[247] +48 * image_in[248] +30 * image_in[249] -7 * image_in[250] -1 * image_in[251] -5 * image_in[252] -7 * image_in[253] +21 * image_in[254] -23 * image_in[255]
                            -46 * image_in[256] -32 * image_in[257] -12 * image_in[258] -11 * image_in[259] +10 * image_in[260] +8 * image_in[261] +24 * image_in[262] +25 * image_in[263] +14 * image_in[264] +1 * image_in[265] -32 * image_in[266] -42 * image_in[267] -10 * image_in[268] -1 * image_in[269] +2 * image_in[270] -24 * image_in[271] -15 * image_in[272] -21 * image_in[274] +6 * image_in[275] +52 * image_in[276] +31 * image_in[277] +3 * image_in[278] +11 * image_in[279] +11 * image_in[281] +26 * image_in[282] -26 * image_in[283] -21 * image_in[284] -4 * image_in[285] -25 * image_in[286] -8 * image_in[287]
                            +14 * image_in[288] +23 * image_in[289] +24 * image_in[290] +24 * image_in[291] +8 * image_in[292] -17 * image_in[293] -38 * image_in[294] -44 * image_in[295] -37 * image_in[296] -27 * image_in[297] -28 * image_in[298] -36 * image_in[299] -35 * image_in[300] -36 * image_in[301] -37 * image_in[302] -21 * image_in[303] +36 * image_in[304] +39 * image_in[305] +34 * image_in[306] -4 * image_in[307] +17 * image_in[308] +13 * image_in[309] +20 * image_in[310] -42 * image_in[311] -16 * image_in[312] -11 * image_in[313] +10 * image_in[314] +11 * image_in[315] +10 * image_in[316] +8 * image_in[317] +1 * image_in[318] -16 * image_in[319]
                            -13 * image_in[320] -22 * image_in[321] -60 * image_in[322] -72 * image_in[323] -42 * image_in[324] -32 * image_in[325] -30 * image_in[326] -35 * image_in[327] -48 * image_in[328] -46 * image_in[329] -73 * image_in[330] -31 * image_in[331] -9 * image_in[332] -11 * image_in[333] -11 * image_in[334] +14 * image_in[335] +10 * image_in[336] +7 * image_in[337] +9 * image_in[338] -2 * image_in[339] -5 * image_in[340] -8 * image_in[341] +21 * image_in[342] +2 * image_in[343] +8 * image_in[344] -9 * image_in[345] +5 * image_in[346] -5 * image_in[347] -10 * image_in[348] -16 * image_in[349] -52 * image_in[350] -51 * image_in[351]
                            -45 * image_in[352] -27 * image_in[353] -10 * image_in[354] -36 * image_in[355] -33 * image_in[356] -43 * image_in[357] -51 * image_in[358] -34 * image_in[359] -23 * image_in[360] -29 * image_in[361] -30 * image_in[362] +13 * image_in[363] -3 * image_in[364] +4 * image_in[365] +13 * image_in[366] -7 * image_in[367] -15 * image_in[368] +3 * image_in[369] +11 * image_in[370] +2 * image_in[371] +6 * image_in[372] +7 * image_in[373] +15 * image_in[374] +10 * image_in[375] +5 * image_in[376] -22 * image_in[377] -43 * image_in[378] -59 * image_in[379] -52 * image_in[380] -23 * image_in[381] -15 * image_in[382] -7 * image_in[383]
                            -10 * image_in[384] -18 * image_in[385] -8 * image_in[386] -8 * image_in[387] -11 * image_in[388] -28 * image_in[389] -41 * image_in[390] -28 * image_in[391] +2 * image_in[392] +30 * image_in[394] -24 * image_in[395] -15 * image_in[396] +22 * image_in[397] +14 * image_in[398] +32 * image_in[399] +15 * image_in[400] +15 * image_in[401] +22 * image_in[402] +11 * image_in[403] -4 * image_in[404] -20 * image_in[405] -35 * image_in[406] -46 * image_in[407] -25 * image_in[408] -22 * image_in[409] -22 * image_in[410] -12 * image_in[411] +18 * image_in[412] +4 * image_in[413] +15 * image_in[414] +7 * image_in[415]
                            +37 * image_in[416] -16 * image_in[417] -23 * image_in[418] -6 * image_in[419] +6 * image_in[420] -13 * image_in[421] -3 * image_in[422] -14 * image_in[423] -22 * image_in[424] +5 * image_in[425] +23 * image_in[427] +24 * image_in[428] +29 * image_in[429] +34 * image_in[430] +21 * image_in[431] -35 * image_in[433] -55 * image_in[434] -46 * image_in[435] -29 * image_in[436] -17 * image_in[437] +13 * image_in[438] +1 * image_in[439] +9 * image_in[440] +10 * image_in[441] -8 * image_in[442] +6 * image_in[443] +17 * image_in[444] +1 * image_in[445] -45 * image_in[446] +4 * image_in[447]
                            -1 * image_in[448] -2 * image_in[449] -39 * image_in[450] +3 * image_in[451] -33 * image_in[452] -4 * image_in[453] -18 * image_in[454] -4 * image_in[455] +13 * image_in[456] +4 * image_in[457] +17 * image_in[458] +29 * image_in[459] -11 * image_in[460] -35 * image_in[461] -45 * image_in[462] -35 * image_in[463] -16 * image_in[464] +7 * image_in[465] +7 * image_in[466] +19 * image_in[467] +15 * image_in[468] +18 * image_in[469] +5 * image_in[470] -17 * image_in[471] -9 * image_in[472] -15 * image_in[473] -58 * image_in[474] -33 * image_in[475] -8 * image_in[477] -31 * image_in[478] -28 * image_in[479]
                            -40 * image_in[480] +2 * image_in[481] +5 * image_in[482] -20 * image_in[483] -20 * image_in[484] -4 * image_in[485] +26 * image_in[486] +13 * image_in[487] -26 * image_in[488] -50 * image_in[489] -29 * image_in[490] +1 * image_in[491] -2 * image_in[492] +22 * image_in[493] +34 * image_in[494] +12 * image_in[495] +12 * image_in[496] -5 * image_in[497] +7 * image_in[498] -18 * image_in[499] +12 * image_in[500] +13 * image_in[501] -41 * image_in[502] -2 * image_in[503] +3 * image_in[504] -15 * image_in[505] -10 * image_in[506] -44 * image_in[507] -9 * image_in[508] -19 * image_in[509] -11 * image_in[510] -9 * image_in[511]
                            -12 * image_in[512] -11 * image_in[513] +5 * image_in[514] -15 * image_in[515] -22 * image_in[516] -32 * image_in[517] -9 * image_in[518] -3 * image_in[519] +16 * image_in[520] +15 * image_in[521] +9 * image_in[522] +5 * image_in[523] -4 * image_in[524] -2 * image_in[525] -11 * image_in[527] +8 * image_in[528] +13 * image_in[529] -21 * image_in[530] -28 * image_in[531] -13 * image_in[533] +20 * image_in[534] -20 * image_in[535] +8 * image_in[536] -15 * image_in[537] +7 * image_in[538] -2 * image_in[539] -7 * image_in[540] -9 * image_in[541] +11 * image_in[542] +17 * image_in[543]
                            +18 * image_in[544] +15 * image_in[545] +11 * image_in[546] +21 * image_in[547] +13 * image_in[548] +7 * image_in[549] +12 * image_in[550] +3 * image_in[551] +9 * image_in[552] +9 * image_in[553] +2 * image_in[554] -10 * image_in[555] +22 * image_in[556] +10 * image_in[557] -27 * image_in[558] -13 * image_in[559] +4 * image_in[560] +12 * image_in[561] +7 * image_in[562] -13 * image_in[563] +1 * image_in[565] -3 * image_in[566] -4 * image_in[567] +9 * image_in[568] +8 * image_in[569] +26 * image_in[570] +30 * image_in[571] +35 * image_in[572] +24 * image_in[573] +22 * image_in[574] +9 * image_in[575]
                            +12 * image_in[576] +9 * image_in[577] +14 * image_in[578] +4 * image_in[579] -4 * image_in[580] +8 * image_in[581] +27 * image_in[582] +15 * image_in[583] -6 * image_in[584] +13 * image_in[585] +33 * image_in[586] +4 * image_in[587] +4 * image_in[588] -4 * image_in[589] -6 * image_in[590] -6 * image_in[591] +7 * image_in[592] -1 * image_in[593] -8 * image_in[594] +9 * image_in[595] +22 * image_in[596] +28 * image_in[597] +29 * image_in[598] +41 * image_in[599] +42 * image_in[600] +32 * image_in[601] +26 * image_in[602] +29 * image_in[603] +14 * image_in[604] +14 * image_in[605] +3 * image_in[606] -5 * image_in[607]
                            +14 * image_in[608] +20 * image_in[609] +33 * image_in[610] +37 * image_in[611] +1 * image_in[612] +4 * image_in[613] +37 * image_in[614] +2 * image_in[615] -3 * image_in[616] +4 * image_in[617] -6 * image_in[618] -16 * image_in[619] +5 * image_in[620] -1 * image_in[621] -3 * image_in[622] -4 * image_in[623] +25 * image_in[624] +21 * image_in[625] +19 * image_in[626] +16 * image_in[627] +36 * image_in[628] +27 * image_in[629] +29 * image_in[630] +15 * image_in[631] +13 * image_in[632] +2 * image_in[633] +10 * image_in[634] +3 * image_in[635] +11 * image_in[636] +25 * image_in[637] +28 * image_in[638] +11 * image_in[639]
                            -23 * image_in[640] -4 * image_in[641] +27 * image_in[642] -2 * image_in[643] +1 * image_in[644] +6 * image_in[645] -15 * image_in[646] -22 * image_in[647] -11 * image_in[648] +27 * image_in[649] +4 * image_in[650] +2 * image_in[651] +15 * image_in[653] +19 * image_in[654] +17 * image_in[655] +16 * image_in[656] +16 * image_in[657] +24 * image_in[658] +16 * image_in[659] +9 * image_in[660] +11 * image_in[661] +3 * image_in[662] -4 * image_in[663] +11 * image_in[664] +12 * image_in[665] +12 * image_in[666] +3 * image_in[667] +5 * image_in[668] +29 * image_in[669] +10 * image_in[670] +3 * image_in[671]
                            -2 * image_in[672] -6 * image_in[674] -28 * image_in[675] -42 * image_in[676] +5 * image_in[677] +3 * image_in[678] -3 * image_in[679] +4 * image_in[680] +12 * image_in[681] +9 * image_in[682] -3 * image_in[683] +14 * image_in[684] +21 * image_in[685] +12 * image_in[686] +24 * image_in[687] -4 * image_in[688] +20 * image_in[689] -19 * image_in[690] -1 * image_in[691] -7 * image_in[692] -19 * image_in[693] +2 * image_in[694] -8 * image_in[695] +20 * image_in[696] +29 * image_in[697] -5 * image_in[698] -3 * image_in[699] -1 * image_in[700] -3 * image_in[702] +14 * image_in[703]
                            +9 * image_in[704] -15 * image_in[705] -11 * image_in[706] -30 * image_in[707] -22 * image_in[708] -21 * image_in[709] -14 * image_in[710] -5 * image_in[711] +7 * image_in[712] +7 * image_in[713] -8 * image_in[714] +13 * image_in[715] +18 * image_in[716] +23 * image_in[717] +12 * image_in[718] +2 * image_in[719] -21 * image_in[720] +2 * image_in[721] +24 * image_in[722] +10 * image_in[723] +11 * image_in[724] +5 * image_in[725] -2 * image_in[726] +2 * image_in[727] -5 * image_in[728] +4 * image_in[729] +5 * image_in[730] +3 * image_in[731] -7 * image_in[732] -23 * image_in[733] -35 * image_in[734] -50 * image_in[735]
                            -34 * image_in[736] +1 * image_in[737] -2 * image_in[738] +21 * image_in[739] +25 * image_in[740] -16 * image_in[742] +30 * image_in[743] +10 * image_in[744] -10 * image_in[745] -22 * image_in[746] +7 * image_in[747] +2 * image_in[748] -4 * image_in[749] +7 * image_in[750] -9 * image_in[751] -3 * image_in[752] -4 * image_in[753] -3 * image_in[754] -4 * image_in[755] +4 * image_in[756] -1 * image_in[757] -5 * image_in[758] -1 * image_in[759] -2 * image_in[760] +17 * image_in[761] +27 * image_in[762] -8 * image_in[763] -1 * image_in[764] +10 * image_in[765] +19 * image_in[766] +17 * image_in[767]
                            +25 * image_in[768] +36 * image_in[769] -6 * image_in[770] +1 * image_in[771] +9 * image_in[772] +14 * image_in[773] -12 * image_in[774] -4 * image_in[775] +4 * image_in[776] -10 * image_in[777] -11 * image_in[778] +5 * image_in[779] +6 * image_in[780] -4 * image_in[782] -4 * image_in[783];
                        if (layer1_out[7] < 0) layer1_out[7] = 0;
                        layer1_out[8] = 34 +1 * image_in[0] +2 * image_in[1] -1 * image_in[2] -6 * image_in[3] -5 * image_in[4] +4 * image_in[5] -6 * image_in[6] -2 * image_in[7] +3 * image_in[8] +2 * image_in[9] +3 * image_in[10] -2 * image_in[11] +7 * image_in[13] -7 * image_in[14] -3 * image_in[15] -1 * image_in[17] -5 * image_in[19] -4 * image_in[20] +5 * image_in[21] -1 * image_in[22] -5 * image_in[23] -3 * image_in[24] +5 * image_in[25] -6 * image_in[27] +3 * image_in[28] -6 * image_in[29] +5 * image_in[30] -1 * image_in[31]
                            -5 * image_in[32] +2 * image_in[33] +11 * image_in[34] +27 * image_in[35] +21 * image_in[36] +13 * image_in[37] +20 * image_in[38] +18 * image_in[39] +25 * image_in[40] +48 * image_in[41] -23 * image_in[42] -26 * image_in[43] -13 * image_in[44] +21 * image_in[45] +33 * image_in[46] +20 * image_in[47] +29 * image_in[48] +17 * image_in[49] +20 * image_in[50] +19 * image_in[51] -2 * image_in[52] +4 * image_in[53] +6 * image_in[54] -1 * image_in[55] +1 * image_in[56] -4 * image_in[57] +4 * image_in[58] -2 * image_in[59] +6 * image_in[60] -3 * image_in[61] +32 * image_in[62] +40 * image_in[63]
                            +45 * image_in[64] +36 * image_in[65] +47 * image_in[66] +32 * image_in[67] +39 * image_in[68] -10 * image_in[69] +25 * image_in[70] +1 * image_in[71] +3 * image_in[72] +5 * image_in[73] +10 * image_in[74] +15 * image_in[75] +47 * image_in[76] +32 * image_in[77] +40 * image_in[78] +28 * image_in[79] +11 * image_in[80] -5 * image_in[81] +1 * image_in[82] -4 * image_in[83] +5 * image_in[84] +1 * image_in[85] +13 * image_in[86] +6 * image_in[88] -15 * image_in[89] +25 * image_in[90] +29 * image_in[91] +2 * image_in[92] +25 * image_in[93] +12 * image_in[94] +33 * image_in[95]
                            +15 * image_in[96] +11 * image_in[97] +8 * image_in[98] +20 * image_in[99] -2 * image_in[100] +7 * image_in[101] +5 * image_in[102] +18 * image_in[103] +11 * image_in[104] +12 * image_in[105] +30 * image_in[106] +17 * image_in[107] +26 * image_in[108] -30 * image_in[109] -4 * image_in[110] -2 * image_in[111] +3 * image_in[112] -20 * image_in[114] +1 * image_in[115] +20 * image_in[116] -10 * image_in[117] -2 * image_in[118] +9 * image_in[119] +4 * image_in[120] +15 * image_in[121] +20 * image_in[122] +13 * image_in[123] +1 * image_in[124] -17 * image_in[125] -10 * image_in[126] -6 * image_in[127]
                            -4 * image_in[128] +16 * image_in[129] -5 * image_in[130] +17 * image_in[131] +16 * image_in[132] +22 * image_in[133] +35 * image_in[134] +16 * image_in[135] -14 * image_in[136] -12 * image_in[137] -23 * image_in[138] +2 * image_in[139] -3 * image_in[140] +4 * image_in[141] +1 * image_in[142] -5 * image_in[143] +7 * image_in[144] -33 * image_in[145] +26 * image_in[146] -12 * image_in[147] +6 * image_in[148] +1 * image_in[149] -35 * image_in[151] -17 * image_in[152] -13 * image_in[153] -6 * image_in[154] -15 * image_in[155] -6 * image_in[156] +10 * image_in[157] +20 * image_in[158] +12 * image_in[159]
                            +17 * image_in[160] +8 * image_in[161] -7 * image_in[162] +9 * image_in[163] +14 * image_in[164] -8 * image_in[165] -3 * image_in[166] -5 * image_in[167] +3 * image_in[168] -1 * image_in[169] -5 * image_in[170] -23 * image_in[171] -1 * image_in[172] +8 * image_in[173] -20 * image_in[174] -6 * image_in[175] -29 * image_in[176] -35 * image_in[177] -57 * image_in[178] -53 * image_in[179] -35 * image_in[180] -29 * image_in[181] -16 * image_in[182] -8 * image_in[183] -2 * image_in[185] -5 * image_in[186] -11 * image_in[187] -7 * image_in[188] -5 * image_in[189] -12 * image_in[190] -1 * image_in[191]
                            -32 * image_in[192] -30 * image_in[193] -11 * image_in[194] +5 * image_in[195] -6 * image_in[196] -23 * image_in[197] +1 * image_in[198] -39 * image_in[199] -1 * image_in[200] -20 * image_in[201] -27 * image_in[202] -36 * image_in[203] -53 * image_in[204] -30 * image_in[205] -49 * image_in[206] -43 * image_in[207] -34 * image_in[208] -20 * image_in[209] -5 * image_in[210] -7 * image_in[211] -3 * image_in[212] -1 * image_in[213] -3 * image_in[214] -15 * image_in[215] -14 * image_in[216] -7 * image_in[217] +3 * image_in[218] -32 * image_in[219] -23 * image_in[220] -18 * image_in[221] +9 * image_in[222] -13 * image_in[223]
                            -1 * image_in[224] -5 * image_in[225] -2 * image_in[226] -36 * image_in[227] -39 * image_in[228] -38 * image_in[229] -60 * image_in[230] -60 * image_in[231] -53 * image_in[232] -32 * image_in[233] -39 * image_in[234] -26 * image_in[235] -28 * image_in[236] -13 * image_in[237] -20 * image_in[238] -1 * image_in[239] -10 * image_in[240] -18 * image_in[241] -26 * image_in[242] -17 * image_in[243] -15 * image_in[244] -10 * image_in[245] -35 * image_in[246] -35 * image_in[247] -48 * image_in[248] -51 * image_in[249] -63 * image_in[250] -22 * image_in[251] -15 * image_in[252] -15 * image_in[253] -30 * image_in[254] -32 * image_in[255]
                            -22 * image_in[256] -55 * image_in[257] -36 * image_in[258] -24 * image_in[259] -41 * image_in[260] -30 * image_in[261] -10 * image_in[262] -19 * image_in[263] -9 * image_in[264] +7 * image_in[265] -2 * image_in[266] -11 * image_in[267] -6 * image_in[268] -22 * image_in[269] -16 * image_in[270] -13 * image_in[271] -8 * image_in[272] -32 * image_in[273] -48 * image_in[274] -39 * image_in[275] -54 * image_in[276] -89 * image_in[277] -45 * image_in[278] +6 * image_in[279] -13 * image_in[280] -4 * image_in[281] -39 * image_in[282] -56 * image_in[283] -38 * image_in[284] -25 * image_in[285] -25 * image_in[286] -29 * image_in[287]
                            -23 * image_in[288] -1 * image_in[289] +9 * image_in[290] +10 * image_in[291] +15 * image_in[292] +4 * image_in[293] -31 * image_in[294] -34 * image_in[295] -48 * image_in[296] -16 * image_in[297] -16 * image_in[298] -3 * image_in[299] -2 * image_in[300] -25 * image_in[301] -27 * image_in[302] -51 * image_in[303] -56 * image_in[304] -91 * image_in[305] -56 * image_in[306] -14 * image_in[307] -4 * image_in[308] -11 * image_in[309] -54 * image_in[310] -45 * image_in[311] -43 * image_in[312] -15 * image_in[313] -9 * image_in[314] -28 * image_in[315] -2 * image_in[316] +16 * image_in[317] +1 * image_in[318] +10 * image_in[319]
                            +8 * image_in[320] -25 * image_in[321] -50 * image_in[322] -55 * image_in[323] -33 * image_in[324] -17 * image_in[325] -14 * image_in[326] +10 * image_in[327] +20 * image_in[328] +23 * image_in[329] -10 * image_in[330] -25 * image_in[331] -59 * image_in[332] -83 * image_in[333] -65 * image_in[334] +19 * image_in[335] +6 * image_in[336] -15 * image_in[337] -45 * image_in[338] -74 * image_in[339] -40 * image_in[340] -17 * image_in[341] +8 * image_in[342] -5 * image_in[343] +9 * image_in[344] +13 * image_in[345] +28 * image_in[346] +32 * image_in[347] +15 * image_in[348] -2 * image_in[349] -31 * image_in[350] -36 * image_in[351]
                            -25 * image_in[352] -8 * image_in[353] -5 * image_in[354] +18 * image_in[355] +12 * image_in[356] +29 * image_in[357] +30 * image_in[358] +35 * image_in[359] -6 * image_in[360] -53 * image_in[361] -69 * image_in[362] +12 * image_in[363] +1 * image_in[364] +4 * image_in[365] -44 * image_in[366] -49 * image_in[367] -19 * image_in[368] +13 * image_in[369] +33 * image_in[370] +22 * image_in[371] +31 * image_in[372] +34 * image_in[373] +48 * image_in[374] +41 * image_in[375] -1 * image_in[376] +10 * image_in[377] -2 * image_in[378] -18 * image_in[379] -6 * image_in[380] -7 * image_in[381] +13 * image_in[382] +10 * image_in[383]
                            +22 * image_in[384] +33 * image_in[385] +30 * image_in[386] +36 * image_in[387] +3 * image_in[388] -33 * image_in[389] -27 * image_in[390] -4 * image_in[391] -1 * image_in[392] -13 * image_in[393] -9 * image_in[394] -17 * image_in[395] -5 * image_in[396] +34 * image_in[397] +25 * image_in[398] +50 * image_in[399] +48 * image_in[400] +57 * image_in[401] +43 * image_in[402] +53 * image_in[403] +27 * image_in[404] +15 * image_in[405] +9 * image_in[406] +1 * image_in[407] +6 * image_in[408] +10 * image_in[409] +19 * image_in[410] +17 * image_in[411] +33 * image_in[412] +25 * image_in[413] +33 * image_in[414] +8 * image_in[415]
                            -2 * image_in[416] -5 * image_in[417] -31 * image_in[418] -1 * image_in[419] -6 * image_in[420] -5 * image_in[421] -17 * image_in[422] +6 * image_in[423] +30 * image_in[425] +31 * image_in[426] +46 * image_in[427] +57 * image_in[428] +43 * image_in[429] +46 * image_in[430] +43 * image_in[431] +37 * image_in[432] +14 * image_in[433] +14 * image_in[434] +20 * image_in[435] +28 * image_in[436] +33 * image_in[437] +29 * image_in[438] +38 * image_in[439] +21 * image_in[440] +16 * image_in[441] +6 * image_in[442] -9 * image_in[443] -3 * image_in[444] +21 * image_in[445] -15 * image_in[446] +12 * image_in[447]
                            -2 * image_in[448] -21 * image_in[450] -14 * image_in[451] -28 * image_in[452] +32 * image_in[453] +38 * image_in[454] +49 * image_in[455] +48 * image_in[456] +45 * image_in[457] +52 * image_in[458] +58 * image_in[459] +23 * image_in[460] +10 * image_in[461] +24 * image_in[462] +38 * image_in[463] +40 * image_in[464] +65 * image_in[465] +48 * image_in[466] +42 * image_in[467] +38 * image_in[468] +40 * image_in[469] +4 * image_in[470] -11 * image_in[471] -11 * image_in[472] +10 * image_in[473] -12 * image_in[474] -1 * image_in[476] -1 * image_in[477] +22 * image_in[478] -21 * image_in[479]
                            -53 * image_in[480] +8 * image_in[481] +11 * image_in[482] +33 * image_in[483] +50 * image_in[484] +40 * image_in[485] +52 * image_in[486] +36 * image_in[487] +9 * image_in[488] +12 * image_in[489] +18 * image_in[490] +48 * image_in[491] +56 * image_in[492] +53 * image_in[493] +49 * image_in[494] +33 * image_in[495] +33 * image_in[496] +11 * image_in[497] +16 * image_in[498] -8 * image_in[499] -10 * image_in[500] +22 * image_in[501] -11 * image_in[502] -5 * image_in[503] -3 * image_in[504] +3 * image_in[506] -28 * image_in[507] -23 * image_in[508] -22 * image_in[509] +12 * image_in[510] +39 * image_in[511]
                            +32 * image_in[512] +39 * image_in[513] +31 * image_in[514] +21 * image_in[515] +13 * image_in[516] +1 * image_in[517] +22 * image_in[518] +36 * image_in[519] +42 * image_in[520] +38 * image_in[521] +31 * image_in[522] +26 * image_in[523] +17 * image_in[524] +18 * image_in[525] -1 * image_in[526] +5 * image_in[527] -10 * image_in[528] +31 * image_in[529] -17 * image_in[530] -5 * image_in[531] -3 * image_in[532] -6 * image_in[533] +7 * image_in[534] -21 * image_in[535] +6 * image_in[536] -21 * image_in[537] +3 * image_in[538] +16 * image_in[539] +11 * image_in[540] +1 * image_in[541] +20 * image_in[542] +20 * image_in[543]
                            +16 * image_in[544] +13 * image_in[545] +28 * image_in[546] +41 * image_in[547] +30 * image_in[548] +30 * image_in[549] +4 * image_in[550] +12 * image_in[551] +7 * image_in[552] +16 * image_in[553] +15 * image_in[554] -11 * image_in[555] -33 * image_in[556] -9 * image_in[557] -18 * image_in[558] +7 * image_in[559] -4 * image_in[560] -6 * image_in[561] +5 * image_in[562] +15 * image_in[563] +10 * image_in[564] -14 * image_in[565] -26 * image_in[566] -11 * image_in[568] -3 * image_in[569] -4 * image_in[570] +15 * image_in[571] +14 * image_in[572] -1 * image_in[573] +17 * image_in[574] +11 * image_in[575] -13 * image_in[577] +5 * image_in[578] -1 * image_in[579] -1 * image_in[580] -9 * image_in[581] -17 * image_in[582] -12 * image_in[583] +7 * image_in[584] -8 * image_in[585] -7 * image_in[586] +5 * image_in[587] -5 * image_in[588] -2 * image_in[589] +29 * image_in[590] +11 * image_in[591] -3 * image_in[592] -17 * image_in[593] -23 * image_in[594] -23 * image_in[595] -24 * image_in[596] -19 * image_in[597] -1 * image_in[598] +7 * image_in[599] +19 * image_in[600] +3 * image_in[601] +1 * image_in[602] -11 * image_in[603] -19 * image_in[604] -19 * image_in[605] -30 * image_in[606] -36 * image_in[607]
                            -18 * image_in[608] -7 * image_in[609] +3 * image_in[611] +4 * image_in[612] -26 * image_in[613] +24 * image_in[614] -4 * image_in[615] -2 * image_in[616] -1 * image_in[617] +13 * image_in[618] +17 * image_in[619] +6 * image_in[620] -16 * image_in[621] -30 * image_in[622] -38 * image_in[623] -19 * image_in[624] -20 * image_in[625] -5 * image_in[627] +6 * image_in[628] -16 * image_in[629] -32 * image_in[630] -31 * image_in[631] -28 * image_in[632] -39 * image_in[633] -45 * image_in[634] -36 * image_in[635] -14 * image_in[636] -18 * image_in[637] -3 * image_in[638] -25 * image_in[639]
                            -19 * image_in[640] -28 * image_in[641] -14 * image_in[642] +6 * image_in[643] +3 * image_in[644] -5 * image_in[645] -8 * image_in[646] -9 * image_in[647] -32 * image_in[648] -19 * image_in[649] -27 * image_in[650] -34 * image_in[651] -19 * image_in[652] -29 * image_in[653] -40 * image_in[654] -44 * image_in[655] -45 * image_in[656] -39 * image_in[657] -31 * image_in[658] -37 * image_in[659] -49 * image_in[660] -42 * image_in[661] -27 * image_in[662] -26 * image_in[663] -27 * image_in[664] -2 * image_in[665] +7 * image_in[666] +5 * image_in[667] -19 * image_in[668] -18 * image_in[669] -21 * image_in[670] +4 * image_in[671]
                            +2 * image_in[672] -6 * image_in[673] -1 * image_in[674] -32 * image_in[675] -12 * image_in[676] -13 * image_in[677] -4 * image_in[678] -10 * image_in[679] -22 * image_in[680] -19 * image_in[681] -30 * image_in[682] -45 * image_in[683] -38 * image_in[684] -58 * image_in[685] -50 * image_in[686] -49 * image_in[687] -37 * image_in[688] -19 * image_in[689] -18 * image_in[690] -9 * image_in[691] +6 * image_in[692] -4 * image_in[693] -9 * image_in[694] +6 * image_in[695] +25 * image_in[697] +4 * image_in[698] +6 * image_in[699] +3 * image_in[700] -4 * image_in[701] -5 * image_in[702] -8 * image_in[703]
                            -8 * image_in[704] +19 * image_in[705] -1 * image_in[706] -1 * image_in[707] -32 * image_in[708] -24 * image_in[709] -30 * image_in[710] -14 * image_in[711] -1 * image_in[712] -2 * image_in[713] -2 * image_in[714] -4 * image_in[715] -1 * image_in[716] -26 * image_in[717] -1 * image_in[718] +14 * image_in[719] +31 * image_in[720] +12 * image_in[721] -19 * image_in[722] +3 * image_in[723] -26 * image_in[724] +2 * image_in[726] +1 * image_in[727] -1 * image_in[728] +4 * image_in[729] +6 * image_in[730] +2 * image_in[731] +29 * image_in[732] +39 * image_in[733] +37 * image_in[734] +21 * image_in[735]
                            +4 * image_in[736] -2 * image_in[737] +6 * image_in[738] +4 * image_in[739] +16 * image_in[740] +12 * image_in[741] +24 * image_in[742] +11 * image_in[743] +14 * image_in[744] -7 * image_in[745] +14 * image_in[746] +16 * image_in[747] +23 * image_in[748] +1 * image_in[749] -12 * image_in[750] +18 * image_in[751] +3 * image_in[752] +4 * image_in[754] +5 * image_in[755] -2 * image_in[756] -5 * image_in[757] +2 * image_in[758] +4 * image_in[759] -4 * image_in[760] -14 * image_in[761] -31 * image_in[762] -19 * image_in[763] -29 * image_in[764] +2 * image_in[765] +4 * image_in[767]
                            -1 * image_in[768] -22 * image_in[769] +1 * image_in[770] -14 * image_in[771] +1 * image_in[772] -13 * image_in[773] +10 * image_in[774] +14 * image_in[775] -11 * image_in[776] -17 * image_in[777] +2 * image_in[778] -5 * image_in[779] -1 * image_in[780] -5 * image_in[781] +3 * image_in[782] +2 * image_in[783];
                        if (layer1_out[8] < 0) layer1_out[8] = 0;
                        layer1_out[9] = 99 -1 * image_in[0] +5 * image_in[1] -4 * image_in[2] +1 * image_in[3] +5 * image_in[4] -3 * image_in[5] +5 * image_in[7] +6 * image_in[8] -5 * image_in[9] +1 * image_in[10] -1 * image_in[11] +4 * image_in[12] +4 * image_in[13] +3 * image_in[14] -4 * image_in[15] +5 * image_in[16] -3 * image_in[17] +2 * image_in[18] -3 * image_in[19] +2 * image_in[20] +2 * image_in[21] +2 * image_in[22] +5 * image_in[23] -3 * image_in[24] +1 * image_in[25] -1 * image_in[26] +3 * image_in[27] -3 * image_in[28] -4 * image_in[29] -2 * image_in[30] -3 * image_in[33] +12 * image_in[34] +16 * image_in[35] +16 * image_in[36] +18 * image_in[37] +21 * image_in[38] +33 * image_in[39] +38 * image_in[40] +52 * image_in[41] +22 * image_in[42] +55 * image_in[43] +28 * image_in[44] +33 * image_in[45] +35 * image_in[46] +36 * image_in[47] +33 * image_in[48] +16 * image_in[49] +14 * image_in[50] +12 * image_in[51] +5 * image_in[52] -6 * image_in[53] +1 * image_in[54] +4 * image_in[55] -5 * image_in[56] -5 * image_in[57] -3 * image_in[58] +2 * image_in[59] +10 * image_in[60] +1 * image_in[61] +13 * image_in[62] +40 * image_in[63]
                            +36 * image_in[64] +2 * image_in[65] +37 * image_in[66] +10 * image_in[67] +15 * image_in[68] +28 * image_in[69] +38 * image_in[70] +46 * image_in[71] +40 * image_in[72] +65 * image_in[73] +63 * image_in[74] +46 * image_in[75] +31 * image_in[76] +20 * image_in[77] +16 * image_in[78] +29 * image_in[79] -10 * image_in[80] -10 * image_in[81] -5 * image_in[82] -2 * image_in[83] +1 * image_in[84] -3 * image_in[85] +16 * image_in[86] +2 * image_in[87] -1 * image_in[88] -1 * image_in[89] +26 * image_in[90] +23 * image_in[91] +29 * image_in[92] +11 * image_in[93] +1 * image_in[94] +20 * image_in[95]
                            +24 * image_in[96] +44 * image_in[97] +50 * image_in[98] +59 * image_in[99] +57 * image_in[100] +52 * image_in[101] +47 * image_in[102] +50 * image_in[103] +49 * image_in[104] +21 * image_in[105] +22 * image_in[106] +16 * image_in[107] +24 * image_in[108] +6 * image_in[109] -4 * image_in[110] +6 * image_in[111] -4 * image_in[112] +5 * image_in[113] +5 * image_in[114] +5 * image_in[115] +10 * image_in[116] -13 * image_in[117] -29 * image_in[118] -14 * image_in[119] -2 * image_in[120] +10 * image_in[121] +10 * image_in[122] +24 * image_in[123] +9 * image_in[124] +15 * image_in[125] +14 * image_in[126] +25 * image_in[127]
                            +16 * image_in[128] +18 * image_in[129] +11 * image_in[130] +13 * image_in[131] -11 * image_in[132] +35 * image_in[133] +5 * image_in[134] +11 * image_in[135] -15 * image_in[136] -1 * image_in[137] +17 * image_in[138] -3 * image_in[139] +6 * image_in[140] -4 * image_in[142] -9 * image_in[143] -40 * image_in[144] -25 * image_in[145] +21 * image_in[146] -7 * image_in[147] +11 * image_in[148] -1 * image_in[149] +22 * image_in[150] -7 * image_in[151] +2 * image_in[152] +14 * image_in[153] +18 * image_in[154] +17 * image_in[155] +6 * image_in[156] +2 * image_in[157] +11 * image_in[158] +4 * image_in[159]
                            +10 * image_in[160] +16 * image_in[161] +5 * image_in[162] -8 * image_in[163] -11 * image_in[164] +35 * image_in[165] +3 * image_in[166] -2 * image_in[167] +1 * image_in[169] +26 * image_in[170] -4 * image_in[171] -3 * image_in[172] -4 * image_in[173] -2 * image_in[174] -6 * image_in[175] -4 * image_in[176] -9 * image_in[177] +4 * image_in[179] +5 * image_in[180] +7 * image_in[181] +8 * image_in[182] +2 * image_in[183] +2 * image_in[184] -1 * image_in[185] +18 * image_in[186] +1 * image_in[187] +10 * image_in[188] +14 * image_in[189] +12 * image_in[190] +4 * image_in[191]
                            +22 * image_in[192] +27 * image_in[193] +6 * image_in[194] -25 * image_in[195] +2 * image_in[196] +4 * image_in[197] -19 * image_in[198] -12 * image_in[199] -27 * image_in[200] -4 * image_in[201] -2 * image_in[202] +15 * image_in[203] -18 * image_in[204] -4 * image_in[205] -10 * image_in[206] +13 * image_in[207] +9 * image_in[208] -2 * image_in[209] +19 * image_in[210] +7 * image_in[211] -4 * image_in[212] -8 * image_in[213] +4 * image_in[215] -3 * image_in[216] -11 * image_in[217] -19 * image_in[218] -10 * image_in[219] +4 * image_in[220] +4 * image_in[221] +2 * image_in[222] -7 * image_in[223]
                            +6 * image_in[224] +32 * image_in[225] -7 * image_in[226] -14 * image_in[227] -42 * image_in[228] -18 * image_in[229] -17 * image_in[230] -9 * image_in[231] -7 * image_in[232] -3 * image_in[233] +1 * image_in[234] -1 * image_in[235] +24 * image_in[236] +19 * image_in[237] +33 * image_in[238] +8 * image_in[239] -7 * image_in[240] -20 * image_in[241] -23 * image_in[242] -24 * image_in[243] -9 * image_in[244] -21 * image_in[245] -37 * image_in[246] -13 * image_in[247] -19 * image_in[248] -7 * image_in[249] -16 * image_in[250] -5 * image_in[251] +19 * image_in[252] +27 * image_in[253] +14 * image_in[254] +8 * image_in[255]
                            +8 * image_in[256] -15 * image_in[257] -7 * image_in[258] +5 * image_in[259] +11 * image_in[260] -1 * image_in[261] +11 * image_in[262] +30 * image_in[263] +41 * image_in[264] +60 * image_in[265] +34 * image_in[266] -10 * image_in[267] -41 * image_in[268] -39 * image_in[269] -32 * image_in[270] -35 * image_in[271] -31 * image_in[272] -24 * image_in[273] -20 * image_in[274] -27 * image_in[275] +25 * image_in[276] +9 * image_in[277] -6 * image_in[278] +3 * image_in[279] +11 * image_in[280] +25 * image_in[281] +24 * image_in[282] +28 * image_in[283] -6 * image_in[284] +15 * image_in[286] +17 * image_in[287]
                            +25 * image_in[288] +25 * image_in[289] +33 * image_in[290] +51 * image_in[291] +55 * image_in[292] +69 * image_in[293] +39 * image_in[294] -22 * image_in[295] -49 * image_in[296] -31 * image_in[297] -14 * image_in[298] -33 * image_in[299] -5 * image_in[300] -9 * image_in[301] -2 * image_in[302] +27 * image_in[303] +57 * image_in[304] +36 * image_in[305] +27 * image_in[306] -12 * image_in[307] +6 * image_in[308] +32 * image_in[309] +50 * image_in[310] +19 * image_in[311] +26 * image_in[312] +4 * image_in[313] +24 * image_in[314] +33 * image_in[315] +36 * image_in[316] +28 * image_in[317] +49 * image_in[318] +49 * image_in[319]
                            +60 * image_in[320] +53 * image_in[321] -2 * image_in[322] -48 * image_in[323] -32 * image_in[324] -5 * image_in[325] -4 * image_in[326] -16 * image_in[327] -10 * image_in[328] -3 * image_in[329] -7 * image_in[330] +24 * image_in[331] +25 * image_in[332] -7 * image_in[333] -8 * image_in[334] +24 * image_in[335] +13 * image_in[336] +21 * image_in[337] +45 * image_in[338] +42 * image_in[339] +7 * image_in[340] +10 * image_in[341] +42 * image_in[342] +36 * image_in[343] +41 * image_in[344] +43 * image_in[345] +45 * image_in[346] +42 * image_in[347] +26 * image_in[348] +3 * image_in[349] -36 * image_in[350] -37 * image_in[351]
                            -18 * image_in[352] +3 * image_in[353] +5 * image_in[354] -26 * image_in[355] -20 * image_in[356] -16 * image_in[357] +12 * image_in[358] +28 * image_in[359] +37 * image_in[360] -15 * image_in[361] -12 * image_in[362] +19 * image_in[363] -2 * image_in[364] +14 * image_in[365] +49 * image_in[366] +26 * image_in[367] +4 * image_in[368] +37 * image_in[369] +54 * image_in[370] +48 * image_in[371] +30 * image_in[372] +36 * image_in[373] +22 * image_in[374] +1 * image_in[375] -13 * image_in[376] -50 * image_in[377] -34 * image_in[378] -36 * image_in[379] -19 * image_in[380] -4 * image_in[381] -19 * image_in[382] -15 * image_in[383]
                            -18 * image_in[384] +10 * image_in[385] +28 * image_in[386] +52 * image_in[387] +35 * image_in[388] -4 * image_in[389] -40 * image_in[390] -22 * image_in[391] +16 * image_in[393] +30 * image_in[394] +19 * image_in[395] -5 * image_in[396] +24 * image_in[397] +36 * image_in[398] +34 * image_in[399] +35 * image_in[400] +14 * image_in[401] +11 * image_in[402] -21 * image_in[403] -36 * image_in[404] -52 * image_in[405] -35 * image_in[406] -15 * image_in[407] -22 * image_in[408] -29 * image_in[409] -26 * image_in[410] -22 * image_in[411] +5 * image_in[412] +26 * image_in[413] +46 * image_in[414] +71 * image_in[415]
                            +71 * image_in[416] -8 * image_in[417] -27 * image_in[418] +5 * image_in[419] -4 * image_in[420] +42 * image_in[422] -15 * image_in[423] +38 * image_in[425] +16 * image_in[426] +31 * image_in[427] +13 * image_in[428] +9 * image_in[429] -19 * image_in[430] -33 * image_in[431] -32 * image_in[432] -32 * image_in[433] -24 * image_in[434] -20 * image_in[435] -33 * image_in[436] -38 * image_in[437] -15 * image_in[438] -14 * image_in[439] +20 * image_in[440] +33 * image_in[441] +27 * image_in[442] +64 * image_in[443] +42 * image_in[444] -2 * image_in[445] -51 * image_in[446] -7 * image_in[447]
                            -1 * image_in[448] +4 * image_in[449] +21 * image_in[450] -20 * image_in[451] -6 * image_in[452] -3 * image_in[453] -13 * image_in[454] -7 * image_in[455] -7 * image_in[457] -21 * image_in[458] -18 * image_in[459] -47 * image_in[460] -36 * image_in[461] -22 * image_in[462] -22 * image_in[463] -38 * image_in[464] -37 * image_in[465] -25 * image_in[466] +4 * image_in[467] +9 * image_in[468] +24 * image_in[469] +22 * image_in[470] +36 * image_in[471] +24 * image_in[472] -42 * image_in[473] -55 * image_in[474] -35 * image_in[475] +3 * image_in[476] +10 * image_in[477] -25 * image_in[478] -17 * image_in[479]
                            -29 * image_in[480] -16 * image_in[481] -15 * image_in[482] -19 * image_in[483] -18 * image_in[484] -26 * image_in[485] -6 * image_in[486] -17 * image_in[487] -52 * image_in[488] -59 * image_in[489] -34 * image_in[490] -22 * image_in[491] -29 * image_in[492] -7 * image_in[493] +3 * image_in[495] +6 * image_in[496] +4 * image_in[497] +22 * image_in[498] +22 * image_in[499] +10 * image_in[500] -33 * image_in[501] -46 * image_in[502] -1 * image_in[503] +3 * image_in[504] +9 * image_in[505] +2 * image_in[507] -17 * image_in[508] -33 * image_in[509] -29 * image_in[510] -13 * image_in[511]
                            -8 * image_in[512] -5 * image_in[513] -14 * image_in[514] -36 * image_in[515] -67 * image_in[516] -69 * image_in[517] -24 * image_in[518] -16 * image_in[519] -23 * image_in[520] -7 * image_in[521] +2 * image_in[522] +16 * image_in[523] +3 * image_in[524] +26 * image_in[525] +29 * image_in[526] +9 * image_in[527] -14 * image_in[528] -22 * image_in[529] -35 * image_in[530] -35 * image_in[531] +2 * image_in[532] +5 * image_in[533] +25 * image_in[534] +8 * image_in[535] -14 * image_in[536] -20 * image_in[537] -12 * image_in[538] -13 * image_in[539] -3 * image_in[540] -8 * image_in[541] -9 * image_in[542] -10 * image_in[543]
                            -6 * image_in[544] -14 * image_in[545] +7 * image_in[546] +9 * image_in[547] +29 * image_in[548] +12 * image_in[549] +21 * image_in[550] +17 * image_in[551] +25 * image_in[552] +5 * image_in[553] +9 * image_in[554] -5 * image_in[555] +19 * image_in[556] -19 * image_in[557] -36 * image_in[558] -10 * image_in[559] -2 * image_in[560] +12 * image_in[561] +15 * image_in[562] -12 * image_in[563] -20 * image_in[564] -26 * image_in[565] -17 * image_in[566] -27 * image_in[567] -5 * image_in[568] +1 * image_in[569] +7 * image_in[570] +14 * image_in[571] +22 * image_in[572] +21 * image_in[573] +33 * image_in[574] +36 * image_in[575]
                            +29 * image_in[576] +29 * image_in[577] +21 * image_in[578] +25 * image_in[579] -1 * image_in[581] +16 * image_in[582] +20 * image_in[583] +1 * image_in[584] -20 * image_in[585] +3 * image_in[587] +1 * image_in[588] +3 * image_in[589] -31 * image_in[590] -12 * image_in[591] -5 * image_in[592] -17 * image_in[593] -24 * image_in[594] -18 * image_in[595] -4 * image_in[596] -11 * image_in[597] +4 * image_in[598] +11 * image_in[599] +29 * image_in[600] +32 * image_in[601] +37 * image_in[602] +49 * image_in[603] +36 * image_in[604] +13 * image_in[605] +24 * image_in[606] +8 * image_in[607] +6 * image_in[609] +7 * image_in[610] -13 * image_in[611] -11 * image_in[612] -3 * image_in[613] +7 * image_in[614] +1 * image_in[615] -5 * image_in[616] +4 * image_in[617] -21 * image_in[618] -23 * image_in[619] -12 * image_in[620] -21 * image_in[621] -30 * image_in[622] -28 * image_in[623] -5 * image_in[624] -8 * image_in[625] +9 * image_in[627] +20 * image_in[628] +21 * image_in[629] +34 * image_in[630] +32 * image_in[631] +37 * image_in[632] +28 * image_in[633] +26 * image_in[634] +15 * image_in[635] +17 * image_in[636] +2 * image_in[637] +16 * image_in[638] -10 * image_in[639]
                            -15 * image_in[640] -5 * image_in[641] +13 * image_in[642] -2 * image_in[643] -5 * image_in[644] +4 * image_in[645] +8 * image_in[647] -37 * image_in[648] -23 * image_in[649] -25 * image_in[650] -10 * image_in[651] -29 * image_in[652] -11 * image_in[653] +13 * image_in[654] +8 * image_in[655] +17 * image_in[656] +8 * image_in[657] +37 * image_in[658] +34 * image_in[659] +14 * image_in[660] +17 * image_in[661] +6 * image_in[662] -10 * image_in[663] -6 * image_in[664] -16 * image_in[665] -16 * image_in[666] -34 * image_in[667] -1 * image_in[668] -12 * image_in[669] +5 * image_in[670] +3 * image_in[671]
                            -2 * image_in[672] +4 * image_in[673] +3 * image_in[674] +18 * image_in[675] -7 * image_in[676] -10 * image_in[677] -15 * image_in[678] +5 * image_in[679] +25 * image_in[680] +18 * image_in[681] +23 * image_in[682] +15 * image_in[683] +15 * image_in[684] +13 * image_in[685] +20 * image_in[686] +21 * image_in[687] +6 * image_in[688] +41 * image_in[689] +3 * image_in[690] -7 * image_in[691] -8 * image_in[692] -10 * image_in[693] +7 * image_in[694] +8 * image_in[695] +22 * image_in[696] -19 * image_in[697] -5 * image_in[698] +1 * image_in[699] -5 * image_in[700] -1 * image_in[701] +3 * image_in[702] +10 * image_in[703]
                            +13 * image_in[704] +10 * image_in[705] +30 * image_in[706] +40 * image_in[707] +67 * image_in[708] +44 * image_in[709] +5 * image_in[710] +15 * image_in[711] +36 * image_in[712] +4 * image_in[713] -6 * image_in[714] +10 * image_in[715] +23 * image_in[716] +31 * image_in[717] +36 * image_in[718] +65 * image_in[719] +16 * image_in[720] +46 * image_in[721] +53 * image_in[722] +45 * image_in[723] +40 * image_in[724] +4 * image_in[725] -1 * image_in[726] -5 * image_in[727] -4 * image_in[729] -2 * image_in[730] +3 * image_in[731] +3 * image_in[732] -21 * image_in[733] +5 * image_in[734] +15 * image_in[735]
                            +52 * image_in[736] +41 * image_in[737] +40 * image_in[738] +62 * image_in[739] +36 * image_in[740] +43 * image_in[741] +32 * image_in[742] +62 * image_in[743] +28 * image_in[744] +46 * image_in[745] +37 * image_in[746] +61 * image_in[747] +28 * image_in[748] +19 * image_in[749] +46 * image_in[750] -8 * image_in[751] -2 * image_in[752] +6 * image_in[753] +4 * image_in[754] +4 * image_in[755] -1 * image_in[756] -3 * image_in[757] +4 * image_in[758] -4 * image_in[759] -2 * image_in[760] +21 * image_in[761] +40 * image_in[762] +17 * image_in[763] +35 * image_in[764] +15 * image_in[765] +27 * image_in[766] +15 * image_in[767]
                            +22 * image_in[768] +61 * image_in[769] +30 * image_in[770] +3 * image_in[771] +11 * image_in[772] +56 * image_in[773] +34 * image_in[774] +19 * image_in[775] +7 * image_in[776] +6 * image_in[777] +24 * image_in[778] +5 * image_in[779] +2 * image_in[780] +5 * image_in[781] +5 * image_in[782] +5 * image_in[783];
                        if (layer1_out[9] < 0) layer1_out[9] = 0;
                        layer1_out[10] = 30 -2 * image_in[0] -4 * image_in[1] -5 * image_in[2] -6 * image_in[3] -2 * image_in[6] +3 * image_in[7] +5 * image_in[8] -4 * image_in[9] -4 * image_in[10] -3 * image_in[11] +1 * image_in[12] +21 * image_in[13] -4 * image_in[14] +5 * image_in[15] -3 * image_in[16] +6 * image_in[17] +3 * image_in[18] -4 * image_in[19] -2 * image_in[20] -4 * image_in[21] +4 * image_in[22] +4 * image_in[23] +3 * image_in[24] -1 * image_in[25] -3 * image_in[26] +1 * image_in[27] -5 * image_in[28] -5 * image_in[29] +5 * image_in[30] -2 * image_in[31]
                            +2 * image_in[32] +3 * image_in[33] -2 * image_in[34] -4 * image_in[35] -9 * image_in[36] +23 * image_in[37] +21 * image_in[38] +21 * image_in[39] +32 * image_in[40] +62 * image_in[41] -9 * image_in[42] -56 * image_in[44] +7 * image_in[45] +26 * image_in[46] +22 * image_in[47] +17 * image_in[48] +22 * image_in[49] +17 * image_in[50] +12 * image_in[51] +2 * image_in[53] +1 * image_in[54] -2 * image_in[55] +5 * image_in[56] -1 * image_in[58] +3 * image_in[59] +16 * image_in[60] -1 * image_in[61] -17 * image_in[62] +1 * image_in[63]
                            -16 * image_in[64] -16 * image_in[65] +4 * image_in[66] -7 * image_in[67] -11 * image_in[68] +17 * image_in[69] +3 * image_in[70] +14 * image_in[71] -11 * image_in[72] +2 * image_in[73] +28 * image_in[74] +27 * image_in[75] +42 * image_in[76] +47 * image_in[77] +25 * image_in[78] +6 * image_in[79] +27 * image_in[80] +18 * image_in[81] -5 * image_in[82] +2 * image_in[83] -5 * image_in[85] +14 * image_in[86] +4 * image_in[87] -2 * image_in[88] +8 * image_in[89] -4 * image_in[90] +1 * image_in[91] -25 * image_in[92] -31 * image_in[93] -15 * image_in[94] -28 * image_in[95]
                            -35 * image_in[96] -23 * image_in[97] -35 * image_in[98] -22 * image_in[99] -10 * image_in[100] -20 * image_in[101] -10 * image_in[102] -18 * image_in[103] -1 * image_in[104] -2 * image_in[105] -6 * image_in[106] +15 * image_in[107] +14 * image_in[108] -17 * image_in[109] -5 * image_in[110] -1 * image_in[111] +4 * image_in[112] +6 * image_in[113] +22 * image_in[114] -5 * image_in[115] +15 * image_in[116] -13 * image_in[117] +5 * image_in[118] -27 * image_in[119] -58 * image_in[120] -58 * image_in[121] -46 * image_in[122] -18 * image_in[123] -18 * image_in[124] +5 * image_in[125] -10 * image_in[126] -8 * image_in[127]
                            -5 * image_in[128] -18 * image_in[129] -1 * image_in[130] +13 * image_in[131] +19 * image_in[132] -1 * image_in[133] -3 * image_in[134] +5 * image_in[135] -32 * image_in[136] -22 * image_in[137] -3 * image_in[138] -2 * image_in[140] +1 * image_in[141] +13 * image_in[143] +1 * image_in[144] +11 * image_in[145] -21 * image_in[146] -32 * image_in[147] -38 * image_in[148] -41 * image_in[149] -47 * image_in[150] -39 * image_in[151] -12 * image_in[152] -5 * image_in[153] -16 * image_in[154] -7 * image_in[155] -31 * image_in[156] -25 * image_in[157] -26 * image_in[158] +11 * image_in[159]
                            -5 * image_in[160] +20 * image_in[161] -9 * image_in[162] -30 * image_in[163] -20 * image_in[164] -40 * image_in[165] -10 * image_in[166] -1 * image_in[167] +3 * image_in[168] +6 * image_in[169] -7 * image_in[170] +25 * image_in[171] -4 * image_in[172] -36 * image_in[173] -7 * image_in[174] -35 * image_in[175] -38 * image_in[176] -47 * image_in[177] -16 * image_in[178] +4 * image_in[179] -1 * image_in[180] +6 * image_in[181] +19 * image_in[182] +14 * image_in[183] +23 * image_in[184] +18 * image_in[185] +30 * image_in[186] +18 * image_in[187] +27 * image_in[188] +16 * image_in[189] +1 * image_in[190] -17 * image_in[191]
                            -35 * image_in[192] -15 * image_in[193] -25 * image_in[194] -7 * image_in[195] -5 * image_in[196] -39 * image_in[197] -8 * image_in[198] +37 * image_in[199] -24 * image_in[200] -45 * image_in[201] -39 * image_in[202] -37 * image_in[203] -51 * image_in[204] -31 * image_in[205] -16 * image_in[206] -11 * image_in[207] +16 * image_in[208] +12 * image_in[209] +29 * image_in[210] +37 * image_in[211] +39 * image_in[212] +31 * image_in[213] +35 * image_in[214] +26 * image_in[215] +30 * image_in[216] +16 * image_in[217] -15 * image_in[218] +7 * image_in[219] -51 * image_in[220] -59 * image_in[221] -34 * image_in[222] +8 * image_in[223] -24 * image_in[225] -24 * image_in[226] -19 * image_in[227] -22 * image_in[228] -39 * image_in[229] -43 * image_in[230] -37 * image_in[231] -39 * image_in[232] -35 * image_in[233] -26 * image_in[234] -13 * image_in[235] +12 * image_in[236] +25 * image_in[237] +38 * image_in[238] +38 * image_in[239] +31 * image_in[240] +21 * image_in[241] +24 * image_in[242] +12 * image_in[243] -12 * image_in[244] +14 * image_in[245] -12 * image_in[246] -26 * image_in[247] -41 * image_in[248] -53 * image_in[249] -5 * image_in[250] -1 * image_in[251] -1 * image_in[252] +1 * image_in[253] -8 * image_in[254] -16 * image_in[255]
                            -37 * image_in[256] -39 * image_in[257] -22 * image_in[258] -33 * image_in[259] -28 * image_in[260] -22 * image_in[261] -12 * image_in[262] -12 * image_in[263] -3 * image_in[264] +24 * image_in[265] +49 * image_in[266] +54 * image_in[267] +23 * image_in[268] +22 * image_in[269] +5 * image_in[270] -5 * image_in[272] -11 * image_in[273] -20 * image_in[274] -53 * image_in[275] -41 * image_in[276] -43 * image_in[277] -5 * image_in[278] +4 * image_in[279] +2 * image_in[280] +21 * image_in[281] +2 * image_in[282] -18 * image_in[283] -16 * image_in[284] -38 * image_in[285] -41 * image_in[286] -38 * image_in[287]
                            -5 * image_in[288] -18 * image_in[289] -15 * image_in[290] -7 * image_in[291] -1 * image_in[292] +34 * image_in[293] +67 * image_in[294] +41 * image_in[295] +25 * image_in[296] +4 * image_in[297] +11 * image_in[298] +5 * image_in[300] -5 * image_in[301] -7 * image_in[302] -3 * image_in[303] -54 * image_in[304] -65 * image_in[305] -31 * image_in[306] +12 * image_in[307] -3 * image_in[308] +10 * image_in[309] +4 * image_in[310] +8 * image_in[311] -6 * image_in[312] -33 * image_in[313] -43 * image_in[314] -18 * image_in[315] +1 * image_in[316] -6 * image_in[317] +8 * image_in[318] +9 * image_in[319]
                            -6 * image_in[320] +61 * image_in[321] +87 * image_in[322] +47 * image_in[323] +30 * image_in[324] +25 * image_in[325] +26 * image_in[326] +12 * image_in[327] +28 * image_in[328] +38 * image_in[329] +19 * image_in[330] +5 * image_in[331] -8 * image_in[332] -30 * image_in[333] +7 * image_in[334] -5 * image_in[336] +7 * image_in[337] +14 * image_in[338] +10 * image_in[339] +20 * image_in[340] +3 * image_in[341] -12 * image_in[342] -11 * image_in[343] +6 * image_in[344] +18 * image_in[345] -13 * image_in[346] -15 * image_in[347] -13 * image_in[348] +55 * image_in[349] +88 * image_in[350] +48 * image_in[351]
                            +25 * image_in[352] +29 * image_in[353] +27 * image_in[354] +23 * image_in[355] +30 * image_in[356] +39 * image_in[357] +34 * image_in[358] +45 * image_in[359] -11 * image_in[360] -39 * image_in[361] -29 * image_in[362] -2 * image_in[363] -1 * image_in[364] -5 * image_in[365] +38 * image_in[366] +32 * image_in[367] +55 * image_in[368] +9 * image_in[369] -10 * image_in[370] +2 * image_in[372] -3 * image_in[373] -16 * image_in[374] -28 * image_in[375] -7 * image_in[376] +38 * image_in[377] +46 * image_in[378] +41 * image_in[379] +17 * image_in[380] +9 * image_in[381] +12 * image_in[382] +19 * image_in[383]
                            +11 * image_in[384] +25 * image_in[385] +4 * image_in[386] -30 * image_in[387] -47 * image_in[388] -72 * image_in[389] -48 * image_in[390] -15 * image_in[391] +6 * image_in[392] +10 * image_in[393] +9 * image_in[394] +37 * image_in[395] +26 * image_in[396] -20 * image_in[397] -21 * image_in[398] -18 * image_in[399] -10 * image_in[400] -18 * image_in[401] -7 * image_in[402] -19 * image_in[403] +4 * image_in[404] +37 * image_in[405] +43 * image_in[406] +32 * image_in[407] +9 * image_in[408] -5 * image_in[409] -2 * image_in[410] -5 * image_in[411] -9 * image_in[412] -11 * image_in[413] -30 * image_in[414] -47 * image_in[415]
                            -82 * image_in[416] -60 * image_in[417] -49 * image_in[418] -6 * image_in[419] -3 * image_in[420] +23 * image_in[421] -19 * image_in[422] -9 * image_in[423] -9 * image_in[424] -13 * image_in[425] -20 * image_in[426] -7 * image_in[427] -12 * image_in[428] -6 * image_in[429] -25 * image_in[430] -14 * image_in[431] +1 * image_in[432] +38 * image_in[433] +36 * image_in[434] +14 * image_in[435] -4 * image_in[436] -18 * image_in[437] +6 * image_in[438] -4 * image_in[439] +12 * image_in[440] -28 * image_in[441] -50 * image_in[442] -67 * image_in[443] -83 * image_in[444] -86 * image_in[445] -45 * image_in[446] -15 * image_in[447]
                            -6 * image_in[448] +4 * image_in[449] +8 * image_in[450] -22 * image_in[451] +12 * image_in[452] -2 * image_in[453] -16 * image_in[454] -19 * image_in[455] +6 * image_in[456] -4 * image_in[457] -8 * image_in[458] +5 * image_in[459] +2 * image_in[460] +21 * image_in[461] +13 * image_in[462] -5 * image_in[463] +4 * image_in[464] -15 * image_in[465] -15 * image_in[466] -4 * image_in[467] -10 * image_in[468] -65 * image_in[469] -75 * image_in[470] -99 * image_in[471] -89 * image_in[472] -97 * image_in[473] -42 * image_in[474] -21 * image_in[475] -5 * image_in[476] +16 * image_in[477] -39 * image_in[478] -32 * image_in[479]
                            -2 * image_in[480] -27 * image_in[481] -45 * image_in[482] -10 * image_in[483] -9 * image_in[484] +8 * image_in[485] +4 * image_in[486] +11 * image_in[487] +14 * image_in[488] +14 * image_in[489] +26 * image_in[490] -6 * image_in[491] -12 * image_in[492] -4 * image_in[493] +7 * image_in[494] +10 * image_in[495] -29 * image_in[496] -35 * image_in[497] -75 * image_in[498] -84 * image_in[499] -73 * image_in[500] -72 * image_in[501] -34 * image_in[502] +6 * image_in[503] -1 * image_in[504] +15 * image_in[505] -7 * image_in[506] -21 * image_in[507] -30 * image_in[508] -49 * image_in[509] -62 * image_in[510] -44 * image_in[511]
                            -19 * image_in[512] -1 * image_in[513] +14 * image_in[515] -1 * image_in[516] +13 * image_in[517] +13 * image_in[518] +6 * image_in[519] -13 * image_in[520] +8 * image_in[521] +33 * image_in[522] +2 * image_in[523] -11 * image_in[524] -46 * image_in[525] -89 * image_in[526] -120 * image_in[527] -95 * image_in[528] -29 * image_in[529] +2 * image_in[530] +2 * image_in[531] +5 * image_in[532] +13 * image_in[533] -23 * image_in[534] -43 * image_in[535] -48 * image_in[536] -36 * image_in[537] -19 * image_in[538] -32 * image_in[539] -28 * image_in[540] -10 * image_in[541] +3 * image_in[542] -5 * image_in[543]
                            +6 * image_in[544] -1 * image_in[545] +17 * image_in[546] +1 * image_in[547] +10 * image_in[548] -1 * image_in[549] +1 * image_in[550] +8 * image_in[551] -28 * image_in[552] -73 * image_in[553] -95 * image_in[554] -103 * image_in[555] -33 * image_in[556] -3 * image_in[557] -7 * image_in[558] -3 * image_in[559] -6 * image_in[560] +4 * image_in[561] -24 * image_in[562] -42 * image_in[563] -37 * image_in[564] -24 * image_in[565] +1 * image_in[567] -4 * image_in[568] -19 * image_in[569] +11 * image_in[570] -13 * image_in[571] +5 * image_in[572] +15 * image_in[573] +9 * image_in[574] -4 * image_in[575]
                            -11 * image_in[576] -9 * image_in[577] -26 * image_in[578] -27 * image_in[579] -57 * image_in[580] -73 * image_in[581] -73 * image_in[582] -68 * image_in[583] -17 * image_in[584] +11 * image_in[585] +1 * image_in[586] -5 * image_in[587] -4 * image_in[588] -37 * image_in[590] -26 * image_in[591] -4 * image_in[592] +6 * image_in[593] +20 * image_in[594] +18 * image_in[595] -2 * image_in[597] +11 * image_in[598] +4 * image_in[599] +2 * image_in[600] +3 * image_in[601] +6 * image_in[602] -3 * image_in[603] -11 * image_in[604] -41 * image_in[605] -47 * image_in[606] -59 * image_in[607]
                            -55 * image_in[608] -55 * image_in[609] -78 * image_in[610] -88 * image_in[611] -10 * image_in[612] +10 * image_in[613] -12 * image_in[614] +2 * image_in[615] +3 * image_in[616] +4 * image_in[617] -45 * image_in[618] -35 * image_in[619] -16 * image_in[620] +48 * image_in[621] +30 * image_in[622] +14 * image_in[623] +7 * image_in[624] +5 * image_in[625] +11 * image_in[626] +4 * image_in[627] +6 * image_in[628] +3 * image_in[629] +11 * image_in[630] -15 * image_in[632] -22 * image_in[633] -53 * image_in[634] -74 * image_in[635] -69 * image_in[636] -55 * image_in[637] -44 * image_in[638] -29 * image_in[639] -9 * image_in[641] +8 * image_in[642] -1 * image_in[643] -4 * image_in[644] +6 * image_in[645] -22 * image_in[646] -43 * image_in[647] -16 * image_in[648] +6 * image_in[649] +17 * image_in[650] +20 * image_in[651] +10 * image_in[652] -2 * image_in[654] +3 * image_in[655] +14 * image_in[656] +29 * image_in[657] +17 * image_in[658] +11 * image_in[659] -6 * image_in[660] -7 * image_in[661] -58 * image_in[662] -67 * image_in[663] -56 * image_in[664] -36 * image_in[665] -26 * image_in[666] -18 * image_in[667] -7 * image_in[668] -16 * image_in[669] +23 * image_in[670] -6 * image_in[671]
                            +4 * image_in[672] -22 * image_in[674] -19 * image_in[675] -16 * image_in[676] +25 * image_in[677] +12 * image_in[678] +4 * image_in[679] +13 * image_in[680] -3 * image_in[681] +14 * image_in[682] +3 * image_in[683] +9 * image_in[684] +7 * image_in[685] +1 * image_in[686] +19 * image_in[687] -9 * image_in[688] -12 * image_in[689] -9 * image_in[690] -12 * image_in[691] -17 * image_in[692] -14 * image_in[693] -3 * image_in[694] +22 * image_in[695] -12 * image_in[696] -28 * image_in[697] +1 * image_in[698] -6 * image_in[699] -4 * image_in[700] +3 * image_in[701] -2 * image_in[702] +5 * image_in[703]
                            +10 * image_in[704] +20 * image_in[705] -2 * image_in[706] +21 * image_in[707] +28 * image_in[708] +28 * image_in[709] -4 * image_in[710] +16 * image_in[711] +15 * image_in[712] +5 * image_in[713] +23 * image_in[714] +12 * image_in[715] +19 * image_in[716] +19 * image_in[717] +36 * image_in[718] +30 * image_in[719] +42 * image_in[720] +52 * image_in[721] +17 * image_in[722] +15 * image_in[723] +23 * image_in[724] -6 * image_in[725] -2 * image_in[726] +4 * image_in[727] +1 * image_in[728] +1 * image_in[729] -3 * image_in[730] +5 * image_in[731] +28 * image_in[732] +33 * image_in[733] +35 * image_in[734] +52 * image_in[735]
                            +65 * image_in[736] +74 * image_in[737] +63 * image_in[738] +67 * image_in[739] +53 * image_in[740] +68 * image_in[741] +94 * image_in[742] +56 * image_in[743] +54 * image_in[744] +74 * image_in[745] +56 * image_in[746] +48 * image_in[747] +48 * image_in[748] +65 * image_in[749] +26 * image_in[750] +8 * image_in[751] -4 * image_in[752] +3 * image_in[753] -1 * image_in[754] +6 * image_in[755] -3 * image_in[756] +1 * image_in[757] -4 * image_in[758] +5 * image_in[759] -1 * image_in[760] -30 * image_in[761] -38 * image_in[762] +14 * image_in[763] +16 * image_in[764] +28 * image_in[765] +24 * image_in[766] +12 * image_in[767]
                            +18 * image_in[768] -1 * image_in[769] +48 * image_in[770] +42 * image_in[771] +36 * image_in[772] +3 * image_in[773] +23 * image_in[774] +16 * image_in[775] +17 * image_in[776] +22 * image_in[777] +13 * image_in[778] -6 * image_in[779] -2 * image_in[780] -6 * image_in[781] -5 * image_in[782];
                        if (layer1_out[10] < 0) layer1_out[10] = 0;
                        layer1_out[11] = 17 -3 * image_in[0] -2 * image_in[1] +5 * image_in[2] +4 * image_in[3] -1 * image_in[4] -2 * image_in[5] -1 * image_in[6] -1 * image_in[7] +5 * image_in[8] -3 * image_in[9] +2 * image_in[10] +6 * image_in[11] -5 * image_in[12] +16 * image_in[13] -5 * image_in[14] -6 * image_in[15] +3 * image_in[16] -6 * image_in[17] -5 * image_in[18] +4 * image_in[19] -5 * image_in[20] -1 * image_in[21] +1 * image_in[22] -3 * image_in[23] +1 * image_in[24] -3 * image_in[25] -3 * image_in[26] +3 * image_in[27] +4 * image_in[28] +5 * image_in[29] +6 * image_in[30] -1 * image_in[31]
                            +2 * image_in[32] -5 * image_in[33] +15 * image_in[34] +30 * image_in[35] +25 * image_in[36] +17 * image_in[37] +16 * image_in[38] +17 * image_in[39] +33 * image_in[40] +41 * image_in[41] -6 * image_in[42] +7 * image_in[43] +29 * image_in[44] +26 * image_in[45] +35 * image_in[46] +20 * image_in[47] +20 * image_in[48] +22 * image_in[49] +24 * image_in[50] +12 * image_in[51] -4 * image_in[52] -5 * image_in[53] +4 * image_in[54] +4 * image_in[55] +2 * image_in[56] -1 * image_in[57] +3 * image_in[58] +3 * image_in[59] +10 * image_in[60] -3 * image_in[61] +30 * image_in[62] +57 * image_in[63]
                            +48 * image_in[64] +57 * image_in[65] +75 * image_in[66] +58 * image_in[67] +62 * image_in[68] +22 * image_in[69] +49 * image_in[70] +14 * image_in[71] +29 * image_in[72] +10 * image_in[73] +21 * image_in[74] +17 * image_in[75] +24 * image_in[76] +4 * image_in[77] +15 * image_in[78] +19 * image_in[79] +10 * image_in[80] +19 * image_in[81] +6 * image_in[82] +4 * image_in[83] -1 * image_in[84] -6 * image_in[85] +7 * image_in[86] +3 * image_in[87] -6 * image_in[88] +24 * image_in[89] +53 * image_in[90] +46 * image_in[91] +13 * image_in[92] +50 * image_in[93] +32 * image_in[94] +32 * image_in[95]
                            +21 * image_in[96] +29 * image_in[97] +10 * image_in[98] +14 * image_in[99] -5 * image_in[100] -4 * image_in[101] -1 * image_in[102] -6 * image_in[103] -3 * image_in[104] -8 * image_in[105] +6 * image_in[106] -3 * image_in[107] +5 * image_in[108] -9 * image_in[109] +6 * image_in[110] -1 * image_in[111] +6 * image_in[112] -2 * image_in[113] -20 * image_in[114] -2 * image_in[115] +4 * image_in[116] +4 * image_in[117] +30 * image_in[118] +13 * image_in[119] +10 * image_in[120] +8 * image_in[121] +27 * image_in[122] +2 * image_in[123] +19 * image_in[124] +11 * image_in[125] -10 * image_in[126] -24 * image_in[127]
                            -33 * image_in[128] -8 * image_in[129] -16 * image_in[130] -32 * image_in[131] -33 * image_in[132] -42 * image_in[133] -38 * image_in[134] -26 * image_in[135] -22 * image_in[136] -11 * image_in[137] -7 * image_in[138] +2 * image_in[139] -2 * image_in[140] +4 * image_in[141] +1 * image_in[142] +38 * image_in[144] +12 * image_in[145] +30 * image_in[146] +23 * image_in[147] +46 * image_in[148] +29 * image_in[149] +26 * image_in[150] +12 * image_in[151] +19 * image_in[152] +7 * image_in[153] +2 * image_in[154] -16 * image_in[155] -7 * image_in[156] -20 * image_in[157] -34 * image_in[158] -41 * image_in[159]
                            -22 * image_in[160] -38 * image_in[161] -39 * image_in[162] -43 * image_in[163] -36 * image_in[164] -6 * image_in[165] -6 * image_in[166] -3 * image_in[167] +2 * image_in[168] -5 * image_in[169] -10 * image_in[170] +4 * image_in[171] +36 * image_in[172] +36 * image_in[173] +48 * image_in[174] +52 * image_in[175] +33 * image_in[176] +52 * image_in[177] +28 * image_in[178] +24 * image_in[179] +21 * image_in[180] +6 * image_in[181] -15 * image_in[182] -5 * image_in[183] -11 * image_in[184] -19 * image_in[185] -33 * image_in[186] -30 * image_in[187] -24 * image_in[188] -7 * image_in[189] -15 * image_in[190] -34 * image_in[191]
                            -28 * image_in[192] +6 * image_in[193] +17 * image_in[194] +16 * image_in[195] -2 * image_in[196] -1 * image_in[197] +46 * image_in[198] +27 * image_in[199] +40 * image_in[200] +45 * image_in[201] +38 * image_in[202] +35 * image_in[203] +29 * image_in[204] +42 * image_in[205] +44 * image_in[206] +39 * image_in[207] +22 * image_in[208] +3 * image_in[209] -15 * image_in[210] -10 * image_in[211] -10 * image_in[212] -10 * image_in[213] -14 * image_in[214] -19 * image_in[215] -5 * image_in[216] +5 * image_in[217] -21 * image_in[218] -27 * image_in[219] +7 * image_in[220] +17 * image_in[221] +27 * image_in[222] +7 * image_in[223]
                            +14 * image_in[224] +24 * image_in[225] +20 * image_in[226] +14 * image_in[227] +50 * image_in[228] +34 * image_in[229] +22 * image_in[230] +30 * image_in[231] +31 * image_in[232] +36 * image_in[233] +36 * image_in[234] +34 * image_in[235] +30 * image_in[236] -4 * image_in[237] +6 * image_in[238] -19 * image_in[240] -18 * image_in[241] -25 * image_in[242] -7 * image_in[243] -3 * image_in[244] -13 * image_in[245] +13 * image_in[246] +6 * image_in[247] -17 * image_in[248] -18 * image_in[249] -22 * image_in[250] -14 * image_in[251] +11 * image_in[252] +36 * image_in[253] +24 * image_in[254] +13 * image_in[255]
                            +45 * image_in[256] +30 * image_in[257] +12 * image_in[258] +19 * image_in[259] +34 * image_in[260] +21 * image_in[261] +8 * image_in[262] +11 * image_in[263] +5 * image_in[264] -7 * image_in[265] +14 * image_in[266] -7 * image_in[267] -16 * image_in[268] -7 * image_in[269] -22 * image_in[270] -10 * image_in[271] +3 * image_in[272] -7 * image_in[273] +5 * image_in[274] +1 * image_in[275] -1 * image_in[276] -31 * image_in[277] +3 * image_in[278] +21 * image_in[279] +11 * image_in[280] +14 * image_in[281] +26 * image_in[282] -3 * image_in[283] +10 * image_in[284] +20 * image_in[285] +19 * image_in[286] +12 * image_in[287]
                            +12 * image_in[288] +17 * image_in[289] +11 * image_in[290] -21 * image_in[291] -33 * image_in[292] -32 * image_in[293] -24 * image_in[294] -18 * image_in[295] -10 * image_in[296] -5 * image_in[297] -5 * image_in[298] -8 * image_in[299] -9 * image_in[300] +1 * image_in[301] +16 * image_in[302] +8 * image_in[303] +15 * image_in[304] -18 * image_in[305] -6 * image_in[306] -16 * image_in[307] +9 * image_in[308] +9 * image_in[309] +11 * image_in[310] -15 * image_in[311] -7 * image_in[312] -7 * image_in[313] -18 * image_in[314] +12 * image_in[315] -12 * image_in[316] -8 * image_in[317] -23 * image_in[318] -28 * image_in[319]
                            -55 * image_in[320] -62 * image_in[321] -42 * image_in[322] -18 * image_in[323] +19 * image_in[324] +1 * image_in[325] -2 * image_in[326] -9 * image_in[327] -15 * image_in[328] -5 * image_in[329] +16 * image_in[330] +26 * image_in[331] +9 * image_in[332] -28 * image_in[333] -60 * image_in[334] +16 * image_in[335] +19 * image_in[336] +1 * image_in[337] +16 * image_in[338] -10 * image_in[339] -27 * image_in[340] -36 * image_in[341] -46 * image_in[342] -29 * image_in[343] -18 * image_in[344] -42 * image_in[345] -50 * image_in[346] -53 * image_in[347] -68 * image_in[348] -80 * image_in[349] -32 * image_in[350] -4 * image_in[351]
                            +16 * image_in[352] +8 * image_in[353] -7 * image_in[354] -19 * image_in[355] -12 * image_in[356] +2 * image_in[357] +6 * image_in[358] +21 * image_in[359] +41 * image_in[360] -15 * image_in[361] -7 * image_in[362] +14 * image_in[363] +5 * image_in[364] +5 * image_in[365] +12 * image_in[366] -18 * image_in[367] -72 * image_in[368] -56 * image_in[369] -67 * image_in[370] -72 * image_in[371] -64 * image_in[372] -64 * image_in[373] -59 * image_in[374] -56 * image_in[375] -63 * image_in[376] -20 * image_in[377] -7 * image_in[378] +16 * image_in[379] +22 * image_in[380] -3 * image_in[381] -21 * image_in[382] -17 * image_in[383]
                            -14 * image_in[384] +11 * image_in[385] +8 * image_in[386] +39 * image_in[387] +58 * image_in[388] +38 * image_in[389] +18 * image_in[390] +31 * image_in[391] +3 * image_in[392] -4 * image_in[393] +11 * image_in[394] -40 * image_in[395] -77 * image_in[396] -57 * image_in[397] -58 * image_in[398] -42 * image_in[399] -62 * image_in[400] -48 * image_in[401] -38 * image_in[402] -15 * image_in[403] -26 * image_in[404] -2 * image_in[405] +18 * image_in[406] +28 * image_in[407] +22 * image_in[408] +6 * image_in[409] +11 * image_in[410] +20 * image_in[411] +12 * image_in[412] +6 * image_in[413] +27 * image_in[414] +41 * image_in[415]
                            +23 * image_in[416] +28 * image_in[417] +35 * image_in[418] -5 * image_in[419] +5 * image_in[420] -24 * image_in[421] -11 * image_in[422] -12 * image_in[423] -70 * image_in[424] -29 * image_in[425] -14 * image_in[426] -32 * image_in[427] -41 * image_in[428] -42 * image_in[429] -22 * image_in[430] +4 * image_in[431] +4 * image_in[432] +28 * image_in[433] +24 * image_in[434] +26 * image_in[435] +10 * image_in[436] +11 * image_in[437] +6 * image_in[438] +9 * image_in[439] +11 * image_in[440] +25 * image_in[441] -1 * image_in[442] +15 * image_in[443] +44 * image_in[444] +49 * image_in[445] +20 * image_in[446] +18 * image_in[447]
                            +2 * image_in[448] -5 * image_in[449] -13 * image_in[450] -12 * image_in[451] -32 * image_in[452] -20 * image_in[453] +5 * image_in[454] -8 * image_in[455] -22 * image_in[456] -17 * image_in[457] -25 * image_in[458] +4 * image_in[459] +34 * image_in[460] +46 * image_in[461] +32 * image_in[462] +27 * image_in[463] +17 * image_in[464] +17 * image_in[465] +9 * image_in[466] +22 * image_in[467] +14 * image_in[468] +23 * image_in[469] +3 * image_in[470] +8 * image_in[471] +39 * image_in[472] +74 * image_in[473] +43 * image_in[474] +25 * image_in[475] -2 * image_in[476] -1 * image_in[477] +6 * image_in[478] -15 * image_in[479]
                            -27 * image_in[480] -6 * image_in[481] +2 * image_in[482] -11 * image_in[483] -25 * image_in[484] -25 * image_in[485] -8 * image_in[486] +33 * image_in[487] +51 * image_in[488] +67 * image_in[489] +30 * image_in[490] +5 * image_in[491] +7 * image_in[492] +14 * image_in[493] +18 * image_in[494] +10 * image_in[495] +4 * image_in[496] -7 * image_in[497] +7 * image_in[498] +14 * image_in[499] +37 * image_in[500] +98 * image_in[501] +41 * image_in[502] -6 * image_in[503] -4 * image_in[504] -7 * image_in[505] -17 * image_in[506] -4 * image_in[507] -14 * image_in[508] -10 * image_in[510] +6 * image_in[511]
                            -29 * image_in[512] -19 * image_in[513] +49 * image_in[515] +76 * image_in[516] +55 * image_in[517] +35 * image_in[518] +26 * image_in[519] +6 * image_in[520] +17 * image_in[521] +17 * image_in[522] +4 * image_in[523] -7 * image_in[524] -20 * image_in[525] -8 * image_in[526] +17 * image_in[527] +49 * image_in[528] +107 * image_in[529] +22 * image_in[530] +16 * image_in[531] -2 * image_in[532] -4 * image_in[533] -22 * image_in[534] -19 * image_in[535] -8 * image_in[536] -18 * image_in[537] -8 * image_in[538] -6 * image_in[539] -22 * image_in[540] -8 * image_in[541] +16 * image_in[542] +46 * image_in[543]
                            +50 * image_in[544] +47 * image_in[545] +42 * image_in[546] +20 * image_in[547] +4 * image_in[548] +3 * image_in[549] -17 * image_in[550] -14 * image_in[551] -13 * image_in[552] -13 * image_in[553] +1 * image_in[554] -3 * image_in[555] +4 * image_in[556] +39 * image_in[557] +23 * image_in[558] +10 * image_in[559] +4 * image_in[560] -22 * image_in[561] -2 * image_in[562] +2 * image_in[563] -5 * image_in[565] -23 * image_in[566] -4 * image_in[567] -8 * image_in[568] -8 * image_in[569] +10 * image_in[570] +22 * image_in[571] +37 * image_in[572] +34 * image_in[573] +26 * image_in[574] +15 * image_in[575]
                            -11 * image_in[576] -12 * image_in[577] -22 * image_in[578] -35 * image_in[579] -39 * image_in[580] -30 * image_in[581] -21 * image_in[582] -17 * image_in[583] +15 * image_in[584] +14 * image_in[585] +10 * image_in[586] -2 * image_in[588] +10 * image_in[589] +4 * image_in[590] +4 * image_in[591] -14 * image_in[592] -32 * image_in[593] -33 * image_in[594] -18 * image_in[595] -5 * image_in[596] +2 * image_in[597] +6 * image_in[598] +7 * image_in[599] +17 * image_in[600] +18 * image_in[601] +28 * image_in[602] +12 * image_in[603] +4 * image_in[604] -36 * image_in[606] -20 * image_in[607]
                            -20 * image_in[608] -26 * image_in[609] -12 * image_in[610] +14 * image_in[611] -10 * image_in[612] -6 * image_in[613] +29 * image_in[614] -5 * image_in[616] +6 * image_in[617] +7 * image_in[618] +6 * image_in[619] +3 * image_in[620] -11 * image_in[622] +2 * image_in[623] +6 * image_in[624] +4 * image_in[625] -6 * image_in[626] -6 * image_in[627] +3 * image_in[628] +6 * image_in[629] -1 * image_in[630] -4 * image_in[631] -16 * image_in[632] -24 * image_in[633] -29 * image_in[634] -15 * image_in[635] -16 * image_in[636] -11 * image_in[637] -18 * image_in[638] -34 * image_in[639]
                            -14 * image_in[640] -1 * image_in[641] -7 * image_in[642] -2 * image_in[643] +5 * image_in[644] +3 * image_in[645] -10 * image_in[646] -36 * image_in[647] -6 * image_in[648] +11 * image_in[649] +19 * image_in[650] +21 * image_in[651] -2 * image_in[652] +8 * image_in[653] -3 * image_in[654] +3 * image_in[655] -8 * image_in[656] -5 * image_in[657] -11 * image_in[658] +7 * image_in[659] -22 * image_in[660] -44 * image_in[661] -16 * image_in[662] -20 * image_in[663] -15 * image_in[664] -4 * image_in[665] -17 * image_in[666] -26 * image_in[667] -28 * image_in[668] +12 * image_in[669] -11 * image_in[670] +3 * image_in[671]
                            +3 * image_in[672] -4 * image_in[673] -15 * image_in[674] -11 * image_in[675] -18 * image_in[676] +24 * image_in[677] +1 * image_in[678] +2 * image_in[679] +17 * image_in[680] +10 * image_in[681] -1 * image_in[682] +7 * image_in[683] +21 * image_in[684] +35 * image_in[685] +20 * image_in[686] +18 * image_in[687] -11 * image_in[688] -9 * image_in[689] -47 * image_in[690] -52 * image_in[691] -32 * image_in[692] -24 * image_in[693] -45 * image_in[694] -57 * image_in[695] -7 * image_in[696] +16 * image_in[697] +5 * image_in[698] +2 * image_in[699] +2 * image_in[700] +2 * image_in[701] -3 * image_in[702] +2 * image_in[703]
                            +17 * image_in[704] -17 * image_in[705] -20 * image_in[706] +8 * image_in[707] +6 * image_in[708] +9 * image_in[709] +12 * image_in[710] +29 * image_in[711] +10 * image_in[712] +6 * image_in[713] +12 * image_in[714] +25 * image_in[715] -1 * image_in[716] -11 * image_in[717] -41 * image_in[718] -65 * image_in[719] -55 * image_in[720] -14 * image_in[721] -45 * image_in[722] -61 * image_in[723] -24 * image_in[724] -4 * image_in[725] -3 * image_in[726] -5 * image_in[727] +4 * image_in[728] -2 * image_in[729] -2 * image_in[730] +5 * image_in[731] -15 * image_in[732] -5 * image_in[733] -32 * image_in[734] +1 * image_in[735]
                            -1 * image_in[736] -1 * image_in[737] -7 * image_in[739] -3 * image_in[740] -13 * image_in[741] +11 * image_in[742] +21 * image_in[743] +1 * image_in[744] -3 * image_in[745] +4 * image_in[746] -26 * image_in[747] -29 * image_in[748] -18 * image_in[749] -8 * image_in[750] -13 * image_in[751] +2 * image_in[752] -3 * image_in[753] -5 * image_in[754] -3 * image_in[755] -3 * image_in[757] +1 * image_in[758] +3 * image_in[759] +4 * image_in[760] +19 * image_in[761] +38 * image_in[762] +17 * image_in[763] +13 * image_in[764] +4 * image_in[765] +29 * image_in[766] +18 * image_in[767]
                            +27 * image_in[768] +52 * image_in[769] +8 * image_in[770] +48 * image_in[771] +55 * image_in[772] +43 * image_in[773] +12 * image_in[774] +6 * image_in[775] -13 * image_in[776] -3 * image_in[777] -2 * image_in[778] -5 * image_in[779] +5 * image_in[780] +5 * image_in[781] -6 * image_in[782] -3 * image_in[783];
                        if (layer1_out[11] < 0) layer1_out[11] = 0;
                        layer1_out[12] = 126 +4 * image_in[0] +1 * image_in[1] +4 * image_in[2] -2 * image_in[3] +1 * image_in[4] +2 * image_in[5] +5 * image_in[6] -5 * image_in[7] +3 * image_in[8] +1 * image_in[9] +4 * image_in[10] +4 * image_in[11] +1 * image_in[13] -3 * image_in[14] -3 * image_in[15] +1 * image_in[16] -4 * image_in[17] +3 * image_in[18] -1 * image_in[19] -1 * image_in[20] +6 * image_in[21] -3 * image_in[22] +6 * image_in[23] -4 * image_in[24] +6 * image_in[25] -5 * image_in[26] -5 * image_in[27] +1 * image_in[28] -1 * image_in[29] +5 * image_in[30] -1 * image_in[31]
                            +3 * image_in[32] +3 * image_in[33] +14 * image_in[34] +32 * image_in[35] +18 * image_in[36] +12 * image_in[37] +14 * image_in[38] -17 * image_in[39] -1 * image_in[40] +3 * image_in[41] +24 * image_in[42] +24 * image_in[43] +5 * image_in[44] +16 * image_in[45] -17 * image_in[46] -3 * image_in[47] +10 * image_in[48] +22 * image_in[49] +22 * image_in[50] +13 * image_in[51] -2 * image_in[52] -1 * image_in[53] +2 * image_in[54] -3 * image_in[55] +1 * image_in[56] +5 * image_in[57] +4 * image_in[58] -6 * image_in[59] +2 * image_in[60] -1 * image_in[61] +21 * image_in[62] +19 * image_in[63]
                            +34 * image_in[64] +15 * image_in[65] +38 * image_in[66] +13 * image_in[67] +18 * image_in[68] +40 * image_in[69] +33 * image_in[70] +39 * image_in[71] +37 * image_in[72] +44 * image_in[73] +7 * image_in[74] +8 * image_in[75] +2 * image_in[76] +3 * image_in[77] -2 * image_in[78] +10 * image_in[79] +10 * image_in[81] -2 * image_in[82] -6 * image_in[83] -6 * image_in[84] -1 * image_in[85] -1 * image_in[86] -4 * image_in[87] +4 * image_in[88] +7 * image_in[89] +26 * image_in[90] +31 * image_in[91] -13 * image_in[92] +5 * image_in[93] -31 * image_in[95]
                            -21 * image_in[96] -28 * image_in[98] -11 * image_in[99] -4 * image_in[100] -32 * image_in[101] -4 * image_in[102] +14 * image_in[103] +6 * image_in[104] +12 * image_in[105] +10 * image_in[106] -5 * image_in[107] -10 * image_in[108] +32 * image_in[109] +5 * image_in[110] +6 * image_in[111] +2 * image_in[112] -4 * image_in[113] +20 * image_in[114] -5 * image_in[115] -3 * image_in[116] +2 * image_in[117] +5 * image_in[118] -22 * image_in[119] -32 * image_in[120] -54 * image_in[121] -53 * image_in[122] -34 * image_in[123] -34 * image_in[124] +6 * image_in[125] -1 * image_in[126] -15 * image_in[127]
                            -22 * image_in[128] -17 * image_in[129] -9 * image_in[130] -22 * image_in[131] -13 * image_in[132] -19 * image_in[133] -22 * image_in[134] +13 * image_in[135] +13 * image_in[136] +21 * image_in[137] -4 * image_in[138] +2 * image_in[139] -3 * image_in[140] +3 * image_in[141] -5 * image_in[142] +19 * image_in[143] +8 * image_in[144] +23 * image_in[145] +6 * image_in[146] -5 * image_in[147] -17 * image_in[148] -26 * image_in[149] -26 * image_in[150] -37 * image_in[151] -35 * image_in[152] -42 * image_in[153] -31 * image_in[154] -41 * image_in[155] -38 * image_in[156] -60 * image_in[157] -36 * image_in[158] -48 * image_in[159]
                            -32 * image_in[160] -27 * image_in[161] -20 * image_in[162] -16 * image_in[163] -2 * image_in[164] -11 * image_in[165] +23 * image_in[166] +2 * image_in[167] -3 * image_in[169] +23 * image_in[171] +18 * image_in[172] -3 * image_in[173] +15 * image_in[174] +3 * image_in[175] -9 * image_in[176] +1 * image_in[177] +1 * image_in[178] +3 * image_in[179] -13 * image_in[180] -6 * image_in[181] -3 * image_in[182] -8 * image_in[183] -6 * image_in[184] -6 * image_in[185] +5 * image_in[186] -8 * image_in[187] +1 * image_in[188] +4 * image_in[189] -17 * image_in[190] -32 * image_in[191]
                            -12 * image_in[192] +2 * image_in[193] +8 * image_in[194] +8 * image_in[195] +4 * image_in[196] -23 * image_in[197] +44 * image_in[198] +36 * image_in[199] -15 * image_in[200] -9 * image_in[201] +11 * image_in[202] +14 * image_in[203] +10 * image_in[204] +14 * image_in[205] +20 * image_in[206] +15 * image_in[207] +30 * image_in[208] +20 * image_in[209] +22 * image_in[210] +10 * image_in[211] +17 * image_in[212] +21 * image_in[213] +20 * image_in[214] +14 * image_in[215] +27 * image_in[216] +17 * image_in[217] +17 * image_in[218] -3 * image_in[219] -11 * image_in[220] -19 * image_in[221] -21 * image_in[222] -6 * image_in[223]
                            +12 * image_in[224] +33 * image_in[225] +8 * image_in[226] +17 * image_in[227] +17 * image_in[228] +5 * image_in[229] +12 * image_in[230] +19 * image_in[231] +21 * image_in[232] -5 * image_in[233] +21 * image_in[234] +36 * image_in[235] +27 * image_in[236] +24 * image_in[237] +35 * image_in[238] +17 * image_in[239] +14 * image_in[240] +39 * image_in[241] +25 * image_in[242] +26 * image_in[243] +25 * image_in[244] +20 * image_in[245] +32 * image_in[246] +11 * image_in[247] +4 * image_in[248] +9 * image_in[249] +15 * image_in[250] +11 * image_in[251] +16 * image_in[252] +27 * image_in[253] +14 * image_in[254] +22 * image_in[255]
                            +18 * image_in[256] +9 * image_in[257] +24 * image_in[258] +8 * image_in[259] +12 * image_in[260] +13 * image_in[261] +16 * image_in[262] +48 * image_in[263] +50 * image_in[264] +33 * image_in[265] +53 * image_in[266] +57 * image_in[267] +35 * image_in[268] +20 * image_in[269] +7 * image_in[270] +1 * image_in[271] -2 * image_in[272] +14 * image_in[273] +8 * image_in[274] -15 * image_in[275] +28 * image_in[276] +51 * image_in[277] +5 * image_in[278] +16 * image_in[279] +16 * image_in[280] +23 * image_in[281] +19 * image_in[282] +22 * image_in[283] -2 * image_in[284] +24 * image_in[285] +26 * image_in[286] +14 * image_in[287]
                            +11 * image_in[288] +10 * image_in[289] +31 * image_in[290] +39 * image_in[291] +42 * image_in[292] +45 * image_in[293] +68 * image_in[294] +69 * image_in[295] +45 * image_in[296] +13 * image_in[297] +5 * image_in[298] -5 * image_in[299] -9 * image_in[300] +10 * image_in[301] +3 * image_in[302] +10 * image_in[303] +31 * image_in[304] +81 * image_in[305] +50 * image_in[306] -13 * image_in[307] +11 * image_in[308] +28 * image_in[309] +40 * image_in[310] +19 * image_in[311] +27 * image_in[312] +15 * image_in[313] -1 * image_in[314] +8 * image_in[315] +1 * image_in[316] +5 * image_in[317] +11 * image_in[318] +15 * image_in[319]
                            +3 * image_in[320] +21 * image_in[321] +38 * image_in[322] +31 * image_in[323] +15 * image_in[324] -5 * image_in[325] +5 * image_in[326] -17 * image_in[327] -19 * image_in[328] -14 * image_in[329] -16 * image_in[330] -23 * image_in[331] -31 * image_in[332] -4 * image_in[333] -8 * image_in[334] -3 * image_in[335] +14 * image_in[336] +15 * image_in[337] +20 * image_in[338] +16 * image_in[339] +22 * image_in[340] +10 * image_in[341] -6 * image_in[342] -1 * image_in[343] -2 * image_in[344] -18 * image_in[345] -39 * image_in[346] -50 * image_in[347] -77 * image_in[348] -63 * image_in[349] +12 * image_in[350] +8 * image_in[351]
                            -16 * image_in[352] -26 * image_in[353] -26 * image_in[355] -25 * image_in[356] -37 * image_in[357] -57 * image_in[358] -60 * image_in[359] -56 * image_in[360] +26 * image_in[361] +45 * image_in[362] +5 * image_in[363] -2 * image_in[364] +5 * image_in[365] +30 * image_in[366] +12 * image_in[367] +19 * image_in[368] -10 * image_in[369] -21 * image_in[370] -17 * image_in[371] -24 * image_in[372] -34 * image_in[373] -49 * image_in[374] -82 * image_in[375] -88 * image_in[376] -47 * image_in[377] +12 * image_in[378] +9 * image_in[379] +3 * image_in[380] -3 * image_in[381] +12 * image_in[382] -9 * image_in[383]
                            -15 * image_in[384] -29 * image_in[385] -39 * image_in[386] -49 * image_in[387] -25 * image_in[388] -15 * image_in[389] -8 * image_in[390] +17 * image_in[391] +3 * image_in[392] +12 * image_in[393] +19 * image_in[394] +14 * image_in[395] -15 * image_in[396] -47 * image_in[397] -36 * image_in[398] -36 * image_in[399] -29 * image_in[400] -26 * image_in[401] -27 * image_in[402] -60 * image_in[403] -55 * image_in[404] -19 * image_in[405] +22 * image_in[406] +12 * image_in[407] +10 * image_in[408] +9 * image_in[409] +18 * image_in[410] +19 * image_in[411] +18 * image_in[412] -15 * image_in[413] -8 * image_in[414] -3 * image_in[415]
                            -46 * image_in[416] +4 * image_in[417] +35 * image_in[418] -3 * image_in[419] +4 * image_in[420] -7 * image_in[421] +29 * image_in[422] -4 * image_in[423] -23 * image_in[424] -37 * image_in[425] -10 * image_in[426] -33 * image_in[427] -17 * image_in[428] -30 * image_in[429] -23 * image_in[430] -32 * image_in[431] -32 * image_in[432] -1 * image_in[433] +15 * image_in[434] +10 * image_in[435] +7 * image_in[436] +10 * image_in[437] +25 * image_in[438] -5 * image_in[439] +10 * image_in[440] +21 * image_in[441] -16 * image_in[442] -24 * image_in[443] +6 * image_in[444] +8 * image_in[446] +23 * image_in[447]
                            -3 * image_in[448] +3 * image_in[449] -15 * image_in[450] +2 * image_in[451] +2 * image_in[452] -31 * image_in[453] -10 * image_in[454] -12 * image_in[455] -7 * image_in[456] -12 * image_in[457] -12 * image_in[458] -21 * image_in[459] -21 * image_in[460] +9 * image_in[461] +7 * image_in[462] +5 * image_in[463] +2 * image_in[464] +12 * image_in[465] -1 * image_in[466] +10 * image_in[467] +4 * image_in[468] -3 * image_in[469] -11 * image_in[470] -29 * image_in[471] -16 * image_in[472] +41 * image_in[473] +44 * image_in[474] +27 * image_in[475] +1 * image_in[476] +1 * image_in[477] -20 * image_in[478] -20 * image_in[479]
                            -5 * image_in[480] -20 * image_in[481] +20 * image_in[482] +8 * image_in[483] +1 * image_in[484] -3 * image_in[485] -18 * image_in[486] -6 * image_in[487] -3 * image_in[488] +31 * image_in[489] +23 * image_in[490] +19 * image_in[491] +2 * image_in[493] -9 * image_in[494] -15 * image_in[495] +1 * image_in[496] -14 * image_in[497] -23 * image_in[498] -4 * image_in[499] +8 * image_in[500] +40 * image_in[501] +41 * image_in[502] -4 * image_in[503] -2 * image_in[504] +1 * image_in[505] -17 * image_in[506] -13 * image_in[507] -6 * image_in[508] -4 * image_in[509] +15 * image_in[510] +20 * image_in[511]
                            +10 * image_in[512] +6 * image_in[513] -24 * image_in[514] -9 * image_in[515] +10 * image_in[516] +35 * image_in[517] +35 * image_in[518] +10 * image_in[519] -5 * image_in[520] +4 * image_in[521] -2 * image_in[522] -19 * image_in[523] -20 * image_in[524] -13 * image_in[525] -19 * image_in[526] -1 * image_in[528] +33 * image_in[529] +35 * image_in[530] +11 * image_in[531] -8 * image_in[533] -24 * image_in[535] +12 * image_in[536] -36 * image_in[537] -28 * image_in[538] +11 * image_in[539] +20 * image_in[540] +21 * image_in[541] -13 * image_in[542] +7 * image_in[543]
                            +18 * image_in[544] +27 * image_in[545] +25 * image_in[546] +18 * image_in[547] +3 * image_in[548] -10 * image_in[549] -27 * image_in[550] -15 * image_in[551] -17 * image_in[552] -49 * image_in[553] -19 * image_in[554] +15 * image_in[555] +43 * image_in[556] +68 * image_in[557] +28 * image_in[558] +1 * image_in[559] -1 * image_in[560] -7 * image_in[561] +3 * image_in[562] +1 * image_in[563] -36 * image_in[564] -48 * image_in[565] -45 * image_in[566] -37 * image_in[567] +6 * image_in[569] +10 * image_in[571] +19 * image_in[572] +7 * image_in[573] +19 * image_in[574] -5 * image_in[575]
                            -2 * image_in[576] -10 * image_in[577] -23 * image_in[578] -3 * image_in[579] -25 * image_in[580] -23 * image_in[581] -7 * image_in[582] +14 * image_in[583] +79 * image_in[584] +57 * image_in[585] +26 * image_in[586] +5 * image_in[587] -5 * image_in[588] -6 * image_in[589] +6 * image_in[590] +6 * image_in[591] -8 * image_in[592] -44 * image_in[593] -34 * image_in[594] -32 * image_in[595] +4 * image_in[596] +2 * image_in[597] +21 * image_in[598] +5 * image_in[599] +1 * image_in[600] +3 * image_in[601] -5 * image_in[602] -3 * image_in[603] -3 * image_in[604] -2 * image_in[605] -10 * image_in[606] +9 * image_in[607]
                            +10 * image_in[608] +11 * image_in[609] -25 * image_in[610] -1 * image_in[611] +57 * image_in[612] +58 * image_in[613] -1 * image_in[614] +5 * image_in[616] -1 * image_in[617] -28 * image_in[618] -28 * image_in[619] +18 * image_in[620] +24 * image_in[621] -12 * image_in[622] -6 * image_in[623] +8 * image_in[624] +6 * image_in[625] -11 * image_in[626] -18 * image_in[627] -12 * image_in[628] -27 * image_in[629] -6 * image_in[630] -12 * image_in[631] -1 * image_in[632] -4 * image_in[633] -13 * image_in[634] -1 * image_in[635] +4 * image_in[636] -24 * image_in[637] -19 * image_in[638] -15 * image_in[639]
                            +56 * image_in[640] +26 * image_in[641] +14 * image_in[642] +6 * image_in[643] +4 * image_in[644] -1 * image_in[645] -26 * image_in[646] -58 * image_in[647] +9 * image_in[648] +17 * image_in[649] +20 * image_in[650] +22 * image_in[651] +1 * image_in[652] -6 * image_in[653] -15 * image_in[654] -21 * image_in[655] -18 * image_in[656] -26 * image_in[657] -29 * image_in[658] -10 * image_in[659] -26 * image_in[660] -17 * image_in[661] -19 * image_in[662] -16 * image_in[663] -19 * image_in[664] -43 * image_in[665] +4 * image_in[666] -11 * image_in[667] +31 * image_in[668] +19 * image_in[670] +5 * image_in[671]
                            -2 * image_in[672] +1 * image_in[673] -17 * image_in[674] -6 * image_in[675] +42 * image_in[677] +22 * image_in[678] -1 * image_in[679] +7 * image_in[680] -15 * image_in[681] -25 * image_in[682] -34 * image_in[683] -20 * image_in[684] -24 * image_in[685] -28 * image_in[686] -6 * image_in[687] -30 * image_in[688] +13 * image_in[689] +1 * image_in[691] +14 * image_in[692] +7 * image_in[693] +1 * image_in[694] -8 * image_in[695] +23 * image_in[696] +13 * image_in[697] +5 * image_in[698] +4 * image_in[699] -2 * image_in[700] +4 * image_in[701] -4 * image_in[702] +16 * image_in[703]
                            +21 * image_in[704] +18 * image_in[705] +3 * image_in[706] +11 * image_in[707] +31 * image_in[708] +22 * image_in[709] -6 * image_in[710] +18 * image_in[711] +32 * image_in[712] +15 * image_in[713] +19 * image_in[714] +31 * image_in[715] +30 * image_in[716] +50 * image_in[717] +48 * image_in[718] +52 * image_in[719] +39 * image_in[720] +66 * image_in[721] +24 * image_in[722] +31 * image_in[723] +28 * image_in[724] -5 * image_in[725] -2 * image_in[726] -3 * image_in[727] -5 * image_in[728] -4 * image_in[729] +4 * image_in[730] +1 * image_in[732] +3 * image_in[733] -3 * image_in[734] +19 * image_in[735]
                            +31 * image_in[736] +45 * image_in[737] +38 * image_in[738] +47 * image_in[739] +26 * image_in[740] +60 * image_in[741] +78 * image_in[742] +62 * image_in[743] +52 * image_in[744] +63 * image_in[745] +50 * image_in[746] +52 * image_in[747] +33 * image_in[748] +16 * image_in[749] +48 * image_in[750] +16 * image_in[751] +2 * image_in[752] +1 * image_in[754] -4 * image_in[755] +2 * image_in[756] +4 * image_in[757] -2 * image_in[758] -1 * image_in[759] +3 * image_in[760] +18 * image_in[761] +34 * image_in[762] +27 * image_in[763] +32 * image_in[764] +12 * image_in[765] +50 * image_in[766] +18 * image_in[767]
                            +31 * image_in[768] +44 * image_in[769] +45 * image_in[770] +15 * image_in[771] +10 * image_in[772] +40 * image_in[773] +31 * image_in[774] +12 * image_in[775] +7 * image_in[776] -20 * image_in[777] +6 * image_in[778] -2 * image_in[779] +3 * image_in[780] +6 * image_in[781] -4 * image_in[782] +1 * image_in[783];
                        if (layer1_out[12] < 0) layer1_out[12] = 0;
                        layer1_out[13] = 22 -5 * image_in[0] -4 * image_in[1] +6 * image_in[2] +6 * image_in[3] -2 * image_in[4] +6 * image_in[5] -2 * image_in[6] -4 * image_in[7] -4 * image_in[8] +1 * image_in[10] -4 * image_in[11] +2 * image_in[12] -9 * image_in[13] +1 * image_in[14] -2 * image_in[15] +5 * image_in[16] -3 * image_in[17] +1 * image_in[18] +6 * image_in[19] -1 * image_in[21] -6 * image_in[22] -3 * image_in[23] -6 * image_in[24] +3 * image_in[25] +2 * image_in[26] -3 * image_in[27] -1 * image_in[28] -3 * image_in[29] -1 * image_in[30] -3 * image_in[31]
                            -3 * image_in[32] -2 * image_in[33] -18 * image_in[34] -33 * image_in[35] -33 * image_in[36] -26 * image_in[37] -25 * image_in[38] -37 * image_in[39] -41 * image_in[40] -42 * image_in[41] +2 * image_in[42] -23 * image_in[43] -34 * image_in[44] -25 * image_in[45] -26 * image_in[46] -27 * image_in[47] -20 * image_in[48] -17 * image_in[49] -19 * image_in[50] -19 * image_in[51] +3 * image_in[52] -3 * image_in[53] -6 * image_in[54] -5 * image_in[55] -4 * image_in[56] -3 * image_in[57] +3 * image_in[58] +4 * image_in[59] -16 * image_in[60] +2 * image_in[61] -27 * image_in[62] -36 * image_in[63]
                            -48 * image_in[64] -43 * image_in[65] -59 * image_in[66] -31 * image_in[67] -50 * image_in[68] -23 * image_in[69] -16 * image_in[70] +5 * image_in[71] -21 * image_in[72] -26 * image_in[73] -47 * image_in[74] -13 * image_in[75] +6 * image_in[76] -7 * image_in[77] -20 * image_in[78] -11 * image_in[79] +8 * image_in[80] +8 * image_in[81] -1 * image_in[82] -5 * image_in[84] -5 * image_in[85] -6 * image_in[86] -2 * image_in[87] +2 * image_in[88] -24 * image_in[89] -36 * image_in[90] -39 * image_in[91] -56 * image_in[92] -43 * image_in[93] -43 * image_in[94] -46 * image_in[95]
                            -56 * image_in[96] -47 * image_in[97] -30 * image_in[98] -32 * image_in[99] -14 * image_in[100] -28 * image_in[101] -50 * image_in[102] -44 * image_in[103] -63 * image_in[104] -43 * image_in[105] -35 * image_in[106] -12 * image_in[107] -30 * image_in[108] -18 * image_in[109] -1 * image_in[110] -3 * image_in[111] +2 * image_in[112] -3 * image_in[113] +14 * image_in[114] -4 * image_in[115] +4 * image_in[116] -10 * image_in[117] -9 * image_in[118] -14 * image_in[119] -11 * image_in[120] -19 * image_in[122] -16 * image_in[123] -5 * image_in[124] +20 * image_in[125] +9 * image_in[126] +12 * image_in[127]
                            +30 * image_in[128] +16 * image_in[129] -5 * image_in[130] +24 * image_in[131] +49 * image_in[132] +17 * image_in[133] +19 * image_in[134] -11 * image_in[135] -19 * image_in[136] -19 * image_in[137] -12 * image_in[138] -1 * image_in[139] -5 * image_in[140] +5 * image_in[141] -4 * image_in[142] +2 * image_in[143] +14 * image_in[144] +28 * image_in[145] +5 * image_in[146] +27 * image_in[147] +31 * image_in[148] +23 * image_in[149] +6 * image_in[150] -9 * image_in[151] -4 * image_in[152] -11 * image_in[153] +17 * image_in[154] +18 * image_in[155] +39 * image_in[156] +33 * image_in[157] +35 * image_in[158] +34 * image_in[159]
                            +26 * image_in[160] +24 * image_in[161] +26 * image_in[162] +15 * image_in[163] -6 * image_in[164] -32 * image_in[165] -16 * image_in[166] +4 * image_in[167] -6 * image_in[168] -4 * image_in[169] -7 * image_in[170] +11 * image_in[172] +52 * image_in[173] +46 * image_in[174] +33 * image_in[175] +28 * image_in[176] +11 * image_in[177] -7 * image_in[178] -20 * image_in[179] -31 * image_in[180] -43 * image_in[181] -46 * image_in[182] -41 * image_in[183] -38 * image_in[184] -17 * image_in[185] -26 * image_in[186] -1 * image_in[187] +8 * image_in[188] +26 * image_in[189] +40 * image_in[190] +37 * image_in[191]
                            -21 * image_in[192] -31 * image_in[193] -19 * image_in[194] -15 * image_in[195] +3 * image_in[196] +6 * image_in[197] +48 * image_in[198] +33 * image_in[199] +46 * image_in[200] +44 * image_in[201] +37 * image_in[202] +41 * image_in[203] +5 * image_in[204] -5 * image_in[205] -5 * image_in[206] -31 * image_in[207] -47 * image_in[208] -33 * image_in[209] -61 * image_in[210] -49 * image_in[211] -36 * image_in[212] -28 * image_in[213] -2 * image_in[214] +6 * image_in[215] -4 * image_in[216] +15 * image_in[217] +31 * image_in[218] +23 * image_in[219] -11 * image_in[220] -30 * image_in[221] +3 * image_in[222] +4 * image_in[223]
                            +9 * image_in[224] +16 * image_in[225] +42 * image_in[226] +59 * image_in[227] +66 * image_in[228] +54 * image_in[229] +28 * image_in[230] +36 * image_in[231] -4 * image_in[232] +19 * image_in[233] +1 * image_in[234] +1 * image_in[235] +11 * image_in[236] -7 * image_in[237] -33 * image_in[238] -13 * image_in[239] -20 * image_in[240] +8 * image_in[241] +24 * image_in[242] +10 * image_in[243] +8 * image_in[244] +7 * image_in[246] +13 * image_in[247] -29 * image_in[248] -32 * image_in[249] -24 * image_in[250] -14 * image_in[251] +16 * image_in[252] +24 * image_in[253] +43 * image_in[254] +40 * image_in[255]
                            +36 * image_in[256] +44 * image_in[257] +3 * image_in[258] +2 * image_in[259] -1 * image_in[260] -5 * image_in[261] +7 * image_in[262] +14 * image_in[263] +14 * image_in[264] +21 * image_in[265] -4 * image_in[266] -14 * image_in[267] +18 * image_in[268] +22 * image_in[269] +20 * image_in[270] +10 * image_in[271] +8 * image_in[272] +17 * image_in[273] -2 * image_in[274] -2 * image_in[275] -48 * image_in[276] -74 * image_in[277] -23 * image_in[278] +15 * image_in[279] +19 * image_in[280] +22 * image_in[281] +47 * image_in[282] +12 * image_in[283] +31 * image_in[284] +8 * image_in[285] -16 * image_in[286] -5 * image_in[287]
                            -3 * image_in[288] +11 * image_in[289] +8 * image_in[290] +19 * image_in[291] +27 * image_in[292] +26 * image_in[293] -2 * image_in[294] +13 * image_in[295] +13 * image_in[296] +22 * image_in[297] +15 * image_in[298] +29 * image_in[299] +10 * image_in[300] +19 * image_in[301] +10 * image_in[302] -57 * image_in[303] -85 * image_in[304] -96 * image_in[305] -54 * image_in[306] +16 * image_in[307] +10 * image_in[308] +30 * image_in[309] +54 * image_in[310] +17 * image_in[311] +11 * image_in[312] +5 * image_in[313] +7 * image_in[315] +2 * image_in[316] +19 * image_in[317] +17 * image_in[318] +14 * image_in[319]
                            +36 * image_in[320] -4 * image_in[321] -14 * image_in[322] +6 * image_in[323] +16 * image_in[324] -7 * image_in[325] -2 * image_in[326] +8 * image_in[327] +1 * image_in[328] +9 * image_in[329] +37 * image_in[330] -4 * image_in[331] -24 * image_in[332] -63 * image_in[333] -25 * image_in[334] +10 * image_in[335] +15 * image_in[336] +39 * image_in[337] +41 * image_in[338] +41 * image_in[339] -12 * image_in[340] -17 * image_in[341] -15 * image_in[342] +16 * image_in[343] +26 * image_in[344] +20 * image_in[345] +17 * image_in[346] +21 * image_in[347] +35 * image_in[348] -15 * image_in[349] -26 * image_in[350] -11 * image_in[351]
                            +11 * image_in[352] +3 * image_in[353] +11 * image_in[354] +7 * image_in[355] +13 * image_in[356] +33 * image_in[357] +47 * image_in[358] +31 * image_in[359] +71 * image_in[360] +26 * image_in[361] -21 * image_in[362] -1 * image_in[363] -2 * image_in[364] +19 * image_in[365] +41 * image_in[366] -7 * image_in[367] -38 * image_in[368] -20 * image_in[369] +5 * image_in[370] +10 * image_in[371] +11 * image_in[372] +13 * image_in[373] +14 * image_in[374] +8 * image_in[375] -6 * image_in[376] -34 * image_in[377] -26 * image_in[378] -2 * image_in[379] -3 * image_in[380] +10 * image_in[381] +14 * image_in[382] +8 * image_in[383]
                            +27 * image_in[384] +20 * image_in[385] +25 * image_in[386] +50 * image_in[387] +54 * image_in[388] +66 * image_in[389] +31 * image_in[390] -7 * image_in[391] -4 * image_in[392] +14 * image_in[393] +31 * image_in[394] -18 * image_in[395] -8 * image_in[396] +23 * image_in[397] +10 * image_in[398] +14 * image_in[399] +10 * image_in[400] +3 * image_in[401] +3 * image_in[403] -4 * image_in[404] -20 * image_in[405] +2 * image_in[407] +16 * image_in[408] +20 * image_in[409] +21 * image_in[410] +31 * image_in[411] +11 * image_in[412] +13 * image_in[413] +15 * image_in[414] +29 * image_in[415]
                            +34 * image_in[416] +29 * image_in[417] -7 * image_in[418] -3 * image_in[419] +1 * image_in[420] -13 * image_in[421] +18 * image_in[422] +5 * image_in[423] +5 * image_in[424] +12 * image_in[425] +8 * image_in[426] +13 * image_in[427] +21 * image_in[428] +13 * image_in[429] +4 * image_in[430] -8 * image_in[431] -4 * image_in[432] +5 * image_in[433] +26 * image_in[434] +22 * image_in[435] +15 * image_in[436] +28 * image_in[437] +14 * image_in[438] +24 * image_in[439] +10 * image_in[440] +19 * image_in[441] +31 * image_in[442] +26 * image_in[443] -9 * image_in[444] +9 * image_in[445] +34 * image_in[446] +2 * image_in[447] +1 * image_in[449] -32 * image_in[450] -5 * image_in[451] -13 * image_in[452] -1 * image_in[453] +28 * image_in[454] +47 * image_in[455] +48 * image_in[456] +29 * image_in[457] +12 * image_in[458] -9 * image_in[459] -3 * image_in[460] +20 * image_in[461] +44 * image_in[462] +44 * image_in[463] +22 * image_in[464] +24 * image_in[465] +14 * image_in[466] +13 * image_in[467] +18 * image_in[468] +29 * image_in[469] -7 * image_in[470] +19 * image_in[471] +2 * image_in[472] +28 * image_in[473] +5 * image_in[474] +25 * image_in[475] +3 * image_in[476] -13 * image_in[477] +33 * image_in[478] -20 * image_in[479] -5 * image_in[481] +7 * image_in[482] +24 * image_in[483] +36 * image_in[484] +48 * image_in[485] +24 * image_in[486] +7 * image_in[487] +28 * image_in[488] +39 * image_in[489] +45 * image_in[490] +16 * image_in[491] +25 * image_in[492] +13 * image_in[493] -2 * image_in[494] +2 * image_in[495] +3 * image_in[496] +7 * image_in[497] +4 * image_in[498] -3 * image_in[499] +21 * image_in[500] +26 * image_in[501] -3 * image_in[502] -1 * image_in[504] -5 * image_in[505] -1 * image_in[506] -28 * image_in[507] -9 * image_in[508] -5 * image_in[509] -29 * image_in[510] -1 * image_in[511]
                            +24 * image_in[512] +28 * image_in[513] +8 * image_in[515] +36 * image_in[516] +31 * image_in[517] +31 * image_in[518] +9 * image_in[519] +4 * image_in[520] -7 * image_in[521] -7 * image_in[522] -19 * image_in[523] +2 * image_in[524] -3 * image_in[525] -13 * image_in[526] -6 * image_in[527] -6 * image_in[528] -25 * image_in[529] +18 * image_in[530] +29 * image_in[531] -1 * image_in[532] -9 * image_in[533] +8 * image_in[534] -14 * image_in[535] -3 * image_in[536] -15 * image_in[537] -25 * image_in[538] -19 * image_in[539] -20 * image_in[540] -12 * image_in[541] -3 * image_in[542] +9 * image_in[543]
                            +4 * image_in[544] +8 * image_in[545] +17 * image_in[546] +7 * image_in[547] +3 * image_in[548] -3 * image_in[549] -2 * image_in[550] -18 * image_in[551] -18 * image_in[552] -7 * image_in[553] -16 * image_in[554] -31 * image_in[555] -8 * image_in[556] +45 * image_in[558] +15 * image_in[559] +4 * image_in[560] +10 * image_in[561] +14 * image_in[562] -15 * image_in[563] -14 * image_in[564] -33 * image_in[565] -13 * image_in[566] +1 * image_in[567] -28 * image_in[568] -20 * image_in[569] +9 * image_in[570] +19 * image_in[571] +27 * image_in[572] +13 * image_in[573] +14 * image_in[574] +24 * image_in[575]
                            +2 * image_in[576] +5 * image_in[577] -1 * image_in[578] -6 * image_in[579] -1 * image_in[580] +7 * image_in[581] -25 * image_in[582] -28 * image_in[583] -24 * image_in[584] -35 * image_in[585] +24 * image_in[586] +5 * image_in[587] +3 * image_in[588] +6 * image_in[589] +5 * image_in[590] -13 * image_in[591] -29 * image_in[592] +3 * image_in[593] -20 * image_in[594] -9 * image_in[595] -9 * image_in[596] -2 * image_in[597] -3 * image_in[598] +18 * image_in[599] +15 * image_in[600] +6 * image_in[601] +18 * image_in[602] +16 * image_in[603] +10 * image_in[604] +19 * image_in[605] +8 * image_in[606] +10 * image_in[607]
                            +5 * image_in[608] -2 * image_in[609] -22 * image_in[610] -9 * image_in[611] -30 * image_in[612] -28 * image_in[613] +3 * image_in[614] -2 * image_in[615] +6 * image_in[616] -1 * image_in[617] -6 * image_in[618] -30 * image_in[619] -24 * image_in[620] +35 * image_in[621] +17 * image_in[622] +23 * image_in[623] -6 * image_in[624] -6 * image_in[625] +8 * image_in[626] +1 * image_in[627] +3 * image_in[628] +8 * image_in[629] +13 * image_in[630] +19 * image_in[631] +8 * image_in[632] +16 * image_in[633] +8 * image_in[634] +27 * image_in[635] +1 * image_in[636] +13 * image_in[637] -40 * image_in[638] -31 * image_in[639]
                            -24 * image_in[640] -9 * image_in[641] +21 * image_in[642] -6 * image_in[643] +1 * image_in[644] -3 * image_in[645] -18 * image_in[646] -57 * image_in[647] -23 * image_in[648] -16 * image_in[649] +9 * image_in[650] +8 * image_in[651] -21 * image_in[652] +14 * image_in[653] -2 * image_in[654] +8 * image_in[655] +11 * image_in[656] +22 * image_in[657] +17 * image_in[658] +40 * image_in[659] +42 * image_in[660] +26 * image_in[661] +11 * image_in[662] +10 * image_in[663] +2 * image_in[664] -9 * image_in[665] -42 * image_in[666] -38 * image_in[667] -55 * image_in[668] +4 * image_in[669] +18 * image_in[670] -6 * image_in[671]
                            -2 * image_in[672] +2 * image_in[673] -11 * image_in[674] -36 * image_in[675] -42 * image_in[676] -12 * image_in[677] -26 * image_in[678] -29 * image_in[679] -20 * image_in[680] -12 * image_in[681] -17 * image_in[682] -6 * image_in[683] -2 * image_in[684] -1 * image_in[685] +10 * image_in[686] -1 * image_in[687] +15 * image_in[688] -11 * image_in[689] -1 * image_in[690] -5 * image_in[691] -27 * image_in[692] -28 * image_in[693] -39 * image_in[694] -52 * image_in[695] -29 * image_in[696] +22 * image_in[697] +6 * image_in[698] -5 * image_in[699] -6 * image_in[700] +4 * image_in[701] +3 * image_in[702] +6 * image_in[703] -47 * image_in[705] -34 * image_in[706] -55 * image_in[707] -55 * image_in[708] -48 * image_in[709] -41 * image_in[710] -39 * image_in[711] -55 * image_in[712] -46 * image_in[713] -27 * image_in[714] -21 * image_in[715] -40 * image_in[716] -33 * image_in[717] -34 * image_in[718] -59 * image_in[719] -72 * image_in[720] -68 * image_in[721] -53 * image_in[722] -52 * image_in[723] -42 * image_in[724] -1 * image_in[725] +2 * image_in[726] -3 * image_in[727] +6 * image_in[728] -6 * image_in[729] +2 * image_in[731] -41 * image_in[732] -34 * image_in[733] -46 * image_in[734] -38 * image_in[735]
                            -28 * image_in[736] -46 * image_in[737] -50 * image_in[738] -48 * image_in[739] -71 * image_in[740] -67 * image_in[741] -72 * image_in[742] -56 * image_in[743] -66 * image_in[744] -44 * image_in[745] -57 * image_in[746] -47 * image_in[747] -62 * image_in[748] -65 * image_in[749] -32 * image_in[750] -20 * image_in[751] -5 * image_in[752] -4 * image_in[753] -4 * image_in[754] -4 * image_in[755] +4 * image_in[756] +1 * image_in[757] -5 * image_in[758] +4 * image_in[759] +30 * image_in[761] +39 * image_in[762] -8 * image_in[763] -14 * image_in[764] +1 * image_in[765] -13 * image_in[766] -19 * image_in[767]
                            -12 * image_in[768] +36 * image_in[769] -19 * image_in[770] -11 * image_in[771] +2 * image_in[772] +44 * image_in[773] +10 * image_in[774] -8 * image_in[776] -9 * image_in[777] -12 * image_in[778] +2 * image_in[779] +5 * image_in[780] -4 * image_in[781] +3 * image_in[783];
                        if (layer1_out[13] < 0) layer1_out[13] = 0;
                        layer1_out[14] = -49 -1 * image_in[0] +2 * image_in[1] -3 * image_in[2] -1 * image_in[3] -1 * image_in[4] -1 * image_in[5] +2 * image_in[6] -5 * image_in[7] +6 * image_in[8] -3 * image_in[9] +5 * image_in[10] -2 * image_in[11] -5 * image_in[12] +5 * image_in[13] -2 * image_in[14] -1 * image_in[15] -5 * image_in[16] -1 * image_in[17] +4 * image_in[18] -4 * image_in[19] -6 * image_in[20] -3 * image_in[21] -6 * image_in[22] +3 * image_in[23] +6 * image_in[24] -2 * image_in[25] +1 * image_in[26] +2 * image_in[27] -3 * image_in[28] +1 * image_in[29] -2 * image_in[30] +6 * image_in[31]
                            -1 * image_in[32] +5 * image_in[33] +16 * image_in[34] +30 * image_in[35] +25 * image_in[36] +26 * image_in[37] +26 * image_in[38] +10 * image_in[39] +31 * image_in[40] +54 * image_in[41] -9 * image_in[42] -8 * image_in[43] -41 * image_in[44] +14 * image_in[45] +36 * image_in[46] +26 * image_in[47] +32 * image_in[48] +20 * image_in[49] +16 * image_in[50] +17 * image_in[51] +4 * image_in[52] -6 * image_in[53] -1 * image_in[54] -2 * image_in[55] +5 * image_in[56] -6 * image_in[57] -3 * image_in[58] -5 * image_in[59] +20 * image_in[60] -4 * image_in[61] +32 * image_in[62] +44 * image_in[63]
                            +41 * image_in[64] +12 * image_in[65] +48 * image_in[66] +23 * image_in[67] +34 * image_in[68] +13 * image_in[69] +17 * image_in[70] +18 * image_in[71] +2 * image_in[72] +15 * image_in[73] +28 * image_in[74] +40 * image_in[75] +52 * image_in[76] +37 * image_in[77] +47 * image_in[78] +37 * image_in[79] +1 * image_in[80] -13 * image_in[81] +5 * image_in[83] -4 * image_in[84] +2 * image_in[85] +11 * image_in[86] +2 * image_in[87] -4 * image_in[88] -31 * image_in[89] +24 * image_in[90] +15 * image_in[91] -4 * image_in[92] +30 * image_in[93] +5 * image_in[94] -11 * image_in[95]
                            -3 * image_in[96] +4 * image_in[97] -20 * image_in[98] +4 * image_in[99] -6 * image_in[100] +9 * image_in[101] +25 * image_in[102] +27 * image_in[103] +22 * image_in[104] +50 * image_in[105] +60 * image_in[106] +50 * image_in[107] +41 * image_in[108] -29 * image_in[109] +6 * image_in[111] +6 * image_in[112] +6 * image_in[113] -22 * image_in[114] -5 * image_in[115] +4 * image_in[116] -32 * image_in[117] -8 * image_in[118] -2 * image_in[119] -17 * image_in[120] -3 * image_in[121] -15 * image_in[122] -21 * image_in[123] -11 * image_in[124] -4 * image_in[125] +5 * image_in[126] +10 * image_in[127]
                            +8 * image_in[128] +18 * image_in[129] +13 * image_in[130] +26 * image_in[131] +27 * image_in[132] +31 * image_in[133] +24 * image_in[134] +36 * image_in[135] +10 * image_in[136] -10 * image_in[137] -14 * image_in[138] +3 * image_in[139] +1 * image_in[140] -1 * image_in[141] +3 * image_in[142] -28 * image_in[143] -40 * image_in[144] -53 * image_in[145] -36 * image_in[146] -37 * image_in[147] -14 * image_in[148] -27 * image_in[149] -17 * image_in[150] -23 * image_in[151] -7 * image_in[152] -1 * image_in[153] +13 * image_in[154] -3 * image_in[155] +3 * image_in[156] +13 * image_in[157] +19 * image_in[158] +27 * image_in[159]
                            +28 * image_in[160] +27 * image_in[161] +17 * image_in[162] +26 * image_in[163] +48 * image_in[164] +27 * image_in[165] +22 * image_in[166] -5 * image_in[167] +3 * image_in[168] +3 * image_in[169] +1 * image_in[170] -56 * image_in[171] -45 * image_in[172] -39 * image_in[173] -69 * image_in[174] -23 * image_in[175] -15 * image_in[176] -17 * image_in[177] -26 * image_in[178] -14 * image_in[179] -6 * image_in[180] -8 * image_in[181] -3 * image_in[182] +9 * image_in[183] -10 * image_in[184] +6 * image_in[185] -16 * image_in[186] +6 * image_in[187] +3 * image_in[188] +3 * image_in[189] +5 * image_in[190] +36 * image_in[191]
                            +49 * image_in[192] +66 * image_in[193] +11 * image_in[194] +16 * image_in[195] -3 * image_in[196] -6 * image_in[197] -23 * image_in[198] -53 * image_in[199] -44 * image_in[200] -47 * image_in[201] -52 * image_in[202] -32 * image_in[203] -9 * image_in[204] -14 * image_in[205] +2 * image_in[206] -6 * image_in[207] -5 * image_in[208] -4 * image_in[209] -1 * image_in[210] +5 * image_in[211] -10 * image_in[212] -11 * image_in[213] -6 * image_in[214] -13 * image_in[215] -7 * image_in[216] +6 * image_in[217] +5 * image_in[218] +19 * image_in[219] +44 * image_in[220] +49 * image_in[221] +25 * image_in[222] -1 * image_in[223]
                            -2 * image_in[224] -14 * image_in[225] -30 * image_in[226] -42 * image_in[227] -76 * image_in[228] -42 * image_in[229] -34 * image_in[230] -11 * image_in[231] -1 * image_in[232] +2 * image_in[233] -5 * image_in[234] -7 * image_in[235] +4 * image_in[236] +7 * image_in[237] -9 * image_in[238] -22 * image_in[239] -21 * image_in[240] -30 * image_in[241] -37 * image_in[242] -29 * image_in[243] -39 * image_in[244] +4 * image_in[245] -11 * image_in[246] -8 * image_in[247] +34 * image_in[248] +23 * image_in[249] +18 * image_in[250] +32 * image_in[251] -11 * image_in[252] -18 * image_in[253] -35 * image_in[254] -55 * image_in[255]
                            -70 * image_in[256] -46 * image_in[257] -6 * image_in[258] +6 * image_in[259] +10 * image_in[260] +16 * image_in[261] +3 * image_in[262] +13 * image_in[263] +5 * image_in[264] -27 * image_in[266] -47 * image_in[267] -46 * image_in[268] -48 * image_in[269] -42 * image_in[270] -26 * image_in[271] -25 * image_in[272] -2 * image_in[273] -14 * image_in[274] +21 * image_in[275] +7 * image_in[276] +1 * image_in[278] -15 * image_in[279] -2 * image_in[280] -10 * image_in[281] -35 * image_in[282] -63 * image_in[283] -32 * image_in[284] -46 * image_in[285] -9 * image_in[286] +18 * image_in[287]
                            +32 * image_in[288] +33 * image_in[289] +31 * image_in[290] +28 * image_in[291] +13 * image_in[292] +4 * image_in[293] -37 * image_in[294] -57 * image_in[295] -66 * image_in[296] -52 * image_in[297] -29 * image_in[298] -24 * image_in[299] -20 * image_in[300] +3 * image_in[302] +13 * image_in[303] -1 * image_in[304] -52 * image_in[305] -22 * image_in[306] -22 * image_in[307] +3 * image_in[308] -15 * image_in[309] -50 * image_in[310] -69 * image_in[311] -51 * image_in[312] +25 * image_in[314] +32 * image_in[315] +38 * image_in[316] +46 * image_in[317] +33 * image_in[318] +25 * image_in[319]
                            +34 * image_in[320] +27 * image_in[321] +6 * image_in[322] -36 * image_in[323] -18 * image_in[324] -27 * image_in[325] -18 * image_in[326] -9 * image_in[327] +2 * image_in[328] +18 * image_in[329] +16 * image_in[330] +44 * image_in[331] +48 * image_in[332] -12 * image_in[333] -7 * image_in[334] +16 * image_in[335] -2 * image_in[336] -15 * image_in[337] -33 * image_in[338] -60 * image_in[339] -36 * image_in[340] +3 * image_in[341] +33 * image_in[342] +42 * image_in[343] +34 * image_in[344] +34 * image_in[345] +24 * image_in[346] +26 * image_in[347] +33 * image_in[348] +51 * image_in[349] +4 * image_in[350] -13 * image_in[351] +12 * image_in[353] -3 * image_in[354] -2 * image_in[355] +10 * image_in[356] +47 * image_in[357] +64 * image_in[358] +88 * image_in[359] +56 * image_in[360] -24 * image_in[361] -62 * image_in[362] +15 * image_in[363] -7 * image_in[365] -34 * image_in[366] -52 * image_in[367] -41 * image_in[368] +11 * image_in[369] +33 * image_in[370] +22 * image_in[371] +30 * image_in[372] +20 * image_in[373] +22 * image_in[374] +14 * image_in[375] +30 * image_in[376] +28 * image_in[377] +24 * image_in[378] +34 * image_in[379] +24 * image_in[380] +4 * image_in[381] -2 * image_in[382] +2 * image_in[383]
                            +17 * image_in[384] +43 * image_in[385] +58 * image_in[386] +65 * image_in[387] +24 * image_in[388] -38 * image_in[389] -61 * image_in[390] -33 * image_in[391] +1 * image_in[392] -9 * image_in[393] -8 * image_in[394] -42 * image_in[395] -18 * image_in[396] +11 * image_in[397] +18 * image_in[398] +5 * image_in[399] +7 * image_in[400] +10 * image_in[401] +14 * image_in[402] +28 * image_in[403] +20 * image_in[404] +24 * image_in[405] +19 * image_in[406] +31 * image_in[407] +28 * image_in[408] -1 * image_in[409] -19 * image_in[410] -25 * image_in[411] -21 * image_in[412] +1 * image_in[413] +26 * image_in[414] -1 * image_in[415]
                            -3 * image_in[416] -9 * image_in[417] -45 * image_in[418] +1 * image_in[419] -5 * image_in[420] +2 * image_in[421] -9 * image_in[422] -30 * image_in[423] -60 * image_in[424] -25 * image_in[425] -19 * image_in[426] -2 * image_in[427] +8 * image_in[428] +11 * image_in[429] +5 * image_in[430] +21 * image_in[431] +23 * image_in[432] +41 * image_in[433] +36 * image_in[434] +17 * image_in[435] +17 * image_in[436] -9 * image_in[437] -28 * image_in[438] -31 * image_in[439] -26 * image_in[440] -28 * image_in[441] -29 * image_in[442] -28 * image_in[443] -32 * image_in[444] +2 * image_in[445] -46 * image_in[446] -11 * image_in[447]
                            -1 * image_in[448] +6 * image_in[449] -17 * image_in[450] -18 * image_in[451] -61 * image_in[452] -34 * image_in[453] -8 * image_in[454] +15 * image_in[456] +19 * image_in[457] +20 * image_in[458] +34 * image_in[459] +25 * image_in[460] +15 * image_in[461] +25 * image_in[462] +11 * image_in[463] -3 * image_in[464] -25 * image_in[465] -23 * image_in[466] -40 * image_in[467] -36 * image_in[468] -40 * image_in[469] -34 * image_in[470] -36 * image_in[471] -17 * image_in[472] -18 * image_in[473] -71 * image_in[474] -31 * image_in[475] -1 * image_in[477] -16 * image_in[478] -51 * image_in[479]
                            -88 * image_in[480] -45 * image_in[481] -23 * image_in[482] +12 * image_in[483] +32 * image_in[484] +41 * image_in[485] +50 * image_in[486] +44 * image_in[487] +27 * image_in[488] +19 * image_in[489] +8 * image_in[490] -9 * image_in[491] -8 * image_in[492] -12 * image_in[493] -19 * image_in[494] -22 * image_in[495] -25 * image_in[496] -38 * image_in[497] -10 * image_in[498] -18 * image_in[499] -14 * image_in[500] -36 * image_in[501] -68 * image_in[502] +3 * image_in[503] -4 * image_in[504] -5 * image_in[505] -8 * image_in[506] -37 * image_in[507] -98 * image_in[508] -68 * image_in[509] -28 * image_in[510] +14 * image_in[511]
                            +30 * image_in[512] +45 * image_in[513] +52 * image_in[514] +35 * image_in[515] +44 * image_in[516] +18 * image_in[517] +6 * image_in[518] +4 * image_in[519] -15 * image_in[520] -11 * image_in[521] -20 * image_in[523] -12 * image_in[524] -26 * image_in[525] -24 * image_in[526] -3 * image_in[527] -14 * image_in[528] -24 * image_in[529] -25 * image_in[530] -27 * image_in[531] +1 * image_in[532] -8 * image_in[533] -11 * image_in[534] -66 * image_in[535] -87 * image_in[536] -44 * image_in[537] -10 * image_in[538] +5 * image_in[539] +2 * image_in[540] +42 * image_in[541] +52 * image_in[542] +40 * image_in[543]
                            +25 * image_in[544] +3 * image_in[545] +3 * image_in[546] +9 * image_in[547] +11 * image_in[548] -10 * image_in[549] -3 * image_in[550] -6 * image_in[552] +1 * image_in[553] +7 * image_in[554] +10 * image_in[555] -9 * image_in[556] -51 * image_in[557] -43 * image_in[558] -14 * image_in[559] -4 * image_in[560] -14 * image_in[561] +6 * image_in[562] -51 * image_in[563] -69 * image_in[564] -47 * image_in[565] -36 * image_in[566] +7 * image_in[567] +3 * image_in[568] +24 * image_in[569] +31 * image_in[570] +16 * image_in[571] +15 * image_in[572] +17 * image_in[573] +10 * image_in[574] +20 * image_in[575]
                            +11 * image_in[576] +7 * image_in[577] +11 * image_in[578] +10 * image_in[579] +12 * image_in[580] +14 * image_in[581] +11 * image_in[582] -9 * image_in[583] -38 * image_in[584] -6 * image_in[585] -19 * image_in[586] +1 * image_in[588] +3 * image_in[589] -3 * image_in[590] -26 * image_in[591] -62 * image_in[592] -53 * image_in[593] -33 * image_in[594] -18 * image_in[595] +1 * image_in[596] +16 * image_in[597] +12 * image_in[598] +12 * image_in[599] +35 * image_in[600] +34 * image_in[601] +34 * image_in[602] +21 * image_in[603] +9 * image_in[604] +24 * image_in[605] +16 * image_in[606] +19 * image_in[607]
                            +11 * image_in[608] -4 * image_in[609] +13 * image_in[610] -13 * image_in[611] -19 * image_in[612] -35 * image_in[613] +13 * image_in[614] +1 * image_in[615] +5 * image_in[616] +5 * image_in[617] -22 * image_in[618] -17 * image_in[619] -33 * image_in[620] -41 * image_in[621] -51 * image_in[622] -31 * image_in[623] -19 * image_in[624] -30 * image_in[625] +9 * image_in[626] +6 * image_in[627] +24 * image_in[628] +33 * image_in[629] +30 * image_in[630] +19 * image_in[631] +14 * image_in[632] +11 * image_in[633] +20 * image_in[634] -2 * image_in[635] +1 * image_in[636] -27 * image_in[638] -14 * image_in[639]
                            +11 * image_in[640] +20 * image_in[641] -28 * image_in[642] +3 * image_in[643] +5 * image_in[644] -3 * image_in[645] -3 * image_in[646] -19 * image_in[648] -36 * image_in[649] -58 * image_in[650] -58 * image_in[651] -6 * image_in[652] -19 * image_in[653] -25 * image_in[654] -12 * image_in[655] +8 * image_in[656] +11 * image_in[657] +12 * image_in[658] +12 * image_in[659] +27 * image_in[660] +11 * image_in[661] +13 * image_in[662] +12 * image_in[663] -2 * image_in[664] +6 * image_in[665] -19 * image_in[666] +21 * image_in[667] -5 * image_in[668] +19 * image_in[669] -15 * image_in[670] -1 * image_in[671]
                            -5 * image_in[672] -5 * image_in[673] +5 * image_in[674] -40 * image_in[675] -40 * image_in[676] -40 * image_in[677] -48 * image_in[678] -35 * image_in[679] -5 * image_in[680] +8 * image_in[681] -4 * image_in[682] -4 * image_in[683] +4 * image_in[684] -19 * image_in[685] +6 * image_in[686] +14 * image_in[687] +18 * image_in[688] -2 * image_in[689] +33 * image_in[690] +22 * image_in[691] +12 * image_in[692] +1 * image_in[693] +7 * image_in[694] +31 * image_in[695] -5 * image_in[696] -11 * image_in[697] -4 * image_in[698] +4 * image_in[699] +2 * image_in[700] +1 * image_in[701] +3 * image_in[702] -3 * image_in[703]
                            -23 * image_in[704] -44 * image_in[705] -39 * image_in[706] -7 * image_in[707] -38 * image_in[708] -21 * image_in[709] -3 * image_in[710] -9 * image_in[711] -12 * image_in[712] -5 * image_in[713] +3 * image_in[714] +4 * image_in[715] +23 * image_in[716] +23 * image_in[717] +14 * image_in[718] +4 * image_in[719] +29 * image_in[720] +2 * image_in[721] +14 * image_in[722] +8 * image_in[723] -9 * image_in[724] -6 * image_in[725] -5 * image_in[726] +5 * image_in[727] +2 * image_in[728] +1 * image_in[729] +22 * image_in[732] -7 * image_in[733] -3 * image_in[734] +17 * image_in[735]
                            +22 * image_in[736] -4 * image_in[737] -10 * image_in[738] +1 * image_in[739] +32 * image_in[740] +13 * image_in[741] +17 * image_in[742] +13 * image_in[743] +5 * image_in[744] +5 * image_in[745] +24 * image_in[746] -11 * image_in[747] +3 * image_in[748] -18 * image_in[749] -8 * image_in[750] +8 * image_in[751] -1 * image_in[752] -2 * image_in[753] -1 * image_in[754] -4 * image_in[755] -6 * image_in[756] +1 * image_in[757] +2 * image_in[759] -6 * image_in[760] -9 * image_in[761] -18 * image_in[762] -6 * image_in[763] -29 * image_in[764] +3 * image_in[765] -23 * image_in[766] +10 * image_in[767]
                            +5 * image_in[768] -23 * image_in[769] +6 * image_in[770] +15 * image_in[771] +3 * image_in[772] -15 * image_in[773] -10 * image_in[774] -4 * image_in[775] -7 * image_in[776] -14 * image_in[777] -3 * image_in[779] -2 * image_in[780] +3 * image_in[781] -4 * image_in[782];
                        if (layer1_out[14] < 0) layer1_out[14] = 0;
                        layer1_out[15] = -44 +5 * image_in[0] -2 * image_in[1] -2 * image_in[2] -1 * image_in[3] -3 * image_in[5] -1 * image_in[6] -4 * image_in[7] +5 * image_in[8] -2 * image_in[9] +2 * image_in[10] +3 * image_in[11] +4 * image_in[12] +8 * image_in[13] +2 * image_in[14] +4 * image_in[15] +1 * image_in[16] +2 * image_in[18] -5 * image_in[19] -1 * image_in[21] +6 * image_in[22] +2 * image_in[23] +2 * image_in[24] -4 * image_in[25] +3 * image_in[26] -1 * image_in[27] +3 * image_in[28] -3 * image_in[29] +1 * image_in[30] -3 * image_in[31]
                            -3 * image_in[32] -1 * image_in[33] +12 * image_in[34] +25 * image_in[35] +18 * image_in[36] +8 * image_in[37] +17 * image_in[38] +22 * image_in[39] +35 * image_in[40] +36 * image_in[41] -3 * image_in[42] +9 * image_in[43] +29 * image_in[44] +32 * image_in[45] +10 * image_in[46] +25 * image_in[47] +25 * image_in[48] +3 * image_in[49] +14 * image_in[50] +17 * image_in[51] +1 * image_in[52] -6 * image_in[53] +2 * image_in[54] -3 * image_in[55] -1 * image_in[56] +1 * image_in[57] -3 * image_in[58] -2 * image_in[59] +14 * image_in[60] -3 * image_in[61] +19 * image_in[62] +30 * image_in[63]
                            +38 * image_in[64] +30 * image_in[65] +54 * image_in[66] +33 * image_in[67] +49 * image_in[68] +15 * image_in[69] +11 * image_in[70] +8 * image_in[71] +41 * image_in[72] +56 * image_in[73] +69 * image_in[74] +47 * image_in[75] +19 * image_in[76] +29 * image_in[77] +8 * image_in[78] -5 * image_in[79] -21 * image_in[80] -11 * image_in[81] +1 * image_in[82] +2 * image_in[83] +2 * image_in[84] +4 * image_in[85] +18 * image_in[86] -3 * image_in[87] +1 * image_in[88] +18 * image_in[89] +33 * image_in[90] +40 * image_in[91] +34 * image_in[92] +37 * image_in[93] +48 * image_in[94] +29 * image_in[95]
                            +47 * image_in[96] +40 * image_in[97] +33 * image_in[98] +44 * image_in[99] +32 * image_in[100] +50 * image_in[101] +72 * image_in[102] +62 * image_in[103] +98 * image_in[104] +74 * image_in[105] +59 * image_in[106] +26 * image_in[107] +23 * image_in[108] +20 * image_in[109] +6 * image_in[110] -3 * image_in[111] +2 * image_in[112] -1 * image_in[113] -14 * image_in[114] -1 * image_in[115] +8 * image_in[116] +26 * image_in[117] +4 * image_in[118] +18 * image_in[119] +20 * image_in[120] +24 * image_in[121] +59 * image_in[122] +49 * image_in[123] +43 * image_in[124] +22 * image_in[125] +45 * image_in[126] +30 * image_in[127]
                            +44 * image_in[128] +29 * image_in[129] +59 * image_in[130] +34 * image_in[131] +17 * image_in[132] +30 * image_in[133] +16 * image_in[134] +21 * image_in[135] +49 * image_in[136] +33 * image_in[137] +17 * image_in[138] +5 * image_in[139] +1 * image_in[140] -3 * image_in[141] +5 * image_in[142] -16 * image_in[144] -8 * image_in[145] -1 * image_in[146] +15 * image_in[147] -6 * image_in[148] +11 * image_in[149] +24 * image_in[150] +21 * image_in[151] +19 * image_in[152] +10 * image_in[153] +2 * image_in[154] -1 * image_in[155] +19 * image_in[156] +14 * image_in[157] +5 * image_in[158] +21 * image_in[159]
                            +31 * image_in[160] +23 * image_in[161] +15 * image_in[162] +18 * image_in[163] +31 * image_in[164] +62 * image_in[165] +28 * image_in[166] -6 * image_in[167] +3 * image_in[168] +2 * image_in[169] +8 * image_in[170] +6 * image_in[172] +1 * image_in[174] +17 * image_in[175] +27 * image_in[176] +23 * image_in[177] +10 * image_in[178] +9 * image_in[179] +13 * image_in[180] +13 * image_in[181] +7 * image_in[182] +10 * image_in[183] +6 * image_in[184] -2 * image_in[185] +3 * image_in[186] +9 * image_in[187] +5 * image_in[188] +1 * image_in[190] +17 * image_in[191]
                            +82 * image_in[192] +97 * image_in[193] +39 * image_in[194] +15 * image_in[195] +1 * image_in[196] +34 * image_in[197] -54 * image_in[198] -15 * image_in[199] +22 * image_in[200] +20 * image_in[201] -3 * image_in[202] +19 * image_in[203] +45 * image_in[204] +18 * image_in[205] +10 * image_in[206] -1 * image_in[207] +15 * image_in[208] +1 * image_in[209] +12 * image_in[210] +8 * image_in[211] -4 * image_in[212] -12 * image_in[213] -3 * image_in[214] -6 * image_in[215] -1 * image_in[216] -9 * image_in[217] -7 * image_in[218] +3 * image_in[219] +50 * image_in[220] +71 * image_in[221] +22 * image_in[222] +6 * image_in[223]
                            -14 * image_in[224] -18 * image_in[225] -19 * image_in[226] +3 * image_in[229] +22 * image_in[230] +35 * image_in[231] +10 * image_in[232] +20 * image_in[233] +21 * image_in[234] +13 * image_in[235] +14 * image_in[236] +13 * image_in[237] -2 * image_in[238] -26 * image_in[239] -18 * image_in[240] -23 * image_in[241] -20 * image_in[242] -1 * image_in[243] +8 * image_in[244] +8 * image_in[245] -2 * image_in[246] +2 * image_in[247] +37 * image_in[248] +64 * image_in[249] +70 * image_in[250] +32 * image_in[251] -13 * image_in[252] -14 * image_in[253] -11 * image_in[254] -10 * image_in[255]
                            +12 * image_in[256] +19 * image_in[257] +22 * image_in[258] +23 * image_in[259] +33 * image_in[260] +27 * image_in[261] +3 * image_in[262] +22 * image_in[263] +4 * image_in[264] -4 * image_in[265] +5 * image_in[266] -22 * image_in[267] -45 * image_in[268] -49 * image_in[269] -34 * image_in[270] -20 * image_in[271] +3 * image_in[272] +7 * image_in[273] +20 * image_in[274] +12 * image_in[275] +40 * image_in[276] +101 * image_in[277] +37 * image_in[278] -21 * image_in[279] -8 * image_in[280] -39 * image_in[281] -38 * image_in[282] +37 * image_in[283] +26 * image_in[284] +8 * image_in[285] +18 * image_in[286] +35 * image_in[287]
                            +3 * image_in[288] +10 * image_in[289] +8 * image_in[290] +9 * image_in[291] +10 * image_in[292] +32 * image_in[293] +14 * image_in[294] -18 * image_in[295] -28 * image_in[296] -44 * image_in[297] -33 * image_in[298] -28 * image_in[299] -27 * image_in[300] -19 * image_in[301] -35 * image_in[302] +12 * image_in[303] +43 * image_in[304] +100 * image_in[305] +58 * image_in[306] +9 * image_in[307] -27 * image_in[308] -35 * image_in[309] -25 * image_in[310] -4 * image_in[311] +46 * image_in[312] +16 * image_in[313] +10 * image_in[314] -8 * image_in[315] -5 * image_in[316] -2 * image_in[317] +6 * image_in[318] +17 * image_in[319]
                            +37 * image_in[320] +66 * image_in[321] +56 * image_in[322] -10 * image_in[323] -30 * image_in[324] -24 * image_in[325] -25 * image_in[326] -21 * image_in[327] -42 * image_in[328] -58 * image_in[329] -63 * image_in[330] -40 * image_in[331] +10 * image_in[332] +67 * image_in[333] +55 * image_in[334] +18 * image_in[335] -19 * image_in[336] -14 * image_in[337] -35 * image_in[338] +5 * image_in[339] +22 * image_in[340] +2 * image_in[341] -20 * image_in[342] -12 * image_in[343] -18 * image_in[344] -9 * image_in[345] +18 * image_in[346] +15 * image_in[347] +30 * image_in[348] +41 * image_in[349] +35 * image_in[350] +5 * image_in[351]
                            -12 * image_in[352] -17 * image_in[353] -24 * image_in[354] -20 * image_in[355] -19 * image_in[356] -51 * image_in[357] -83 * image_in[358] -81 * image_in[359] -76 * image_in[360] +7 * image_in[361] +28 * image_in[362] +17 * image_in[363] -1 * image_in[364] -16 * image_in[365] -38 * image_in[366] +2 * image_in[367] -18 * image_in[368] -23 * image_in[369] -39 * image_in[370] -32 * image_in[371] -20 * image_in[372] -7 * image_in[373] -22 * image_in[374] -5 * image_in[375] +26 * image_in[376] +39 * image_in[377] +18 * image_in[378] +5 * image_in[379] -12 * image_in[380] -19 * image_in[381] -4 * image_in[382] -3 * image_in[383]
                            -27 * image_in[384] -51 * image_in[385] -41 * image_in[386] -66 * image_in[387] -53 * image_in[388] -9 * image_in[389] +24 * image_in[390] +17 * image_in[391] -2 * image_in[392] -13 * image_in[393] -28 * image_in[394] +1 * image_in[395] -47 * image_in[396] -54 * image_in[397] -38 * image_in[398] -46 * image_in[399] -26 * image_in[400] -17 * image_in[401] -12 * image_in[402] -17 * image_in[403] +10 * image_in[404] +30 * image_in[405] +24 * image_in[406] +13 * image_in[407] -8 * image_in[408] -14 * image_in[409] -9 * image_in[410] -6 * image_in[411] -11 * image_in[412] -29 * image_in[413] -37 * image_in[414] -41 * image_in[415]
                            -26 * image_in[416] +6 * image_in[417] -4 * image_in[419] +3 * image_in[420] +13 * image_in[421] +15 * image_in[422] -17 * image_in[423] -45 * image_in[424] -71 * image_in[425] -46 * image_in[426] -61 * image_in[427] -48 * image_in[428] -25 * image_in[429] -12 * image_in[430] -10 * image_in[431] +21 * image_in[432] +46 * image_in[433] +38 * image_in[434] +10 * image_in[435] -10 * image_in[436] -15 * image_in[437] -1 * image_in[438] +15 * image_in[439] -11 * image_in[440] -11 * image_in[441] -23 * image_in[442] -10 * image_in[443] +17 * image_in[444] +23 * image_in[445] -19 * image_in[446] +12 * image_in[447]
                            +4 * image_in[448] -6 * image_in[449] +43 * image_in[450] +11 * image_in[451] -11 * image_in[452] -54 * image_in[453] -58 * image_in[454] -76 * image_in[455] -66 * image_in[456] -32 * image_in[457] -25 * image_in[458] -2 * image_in[459] +32 * image_in[460] +36 * image_in[461] +25 * image_in[462] +3 * image_in[463] -10 * image_in[464] +4 * image_in[465] +10 * image_in[466] +27 * image_in[467] -2 * image_in[469] +15 * image_in[470] +32 * image_in[471] +56 * image_in[472] +27 * image_in[473] +9 * image_in[474] -13 * image_in[475] -4 * image_in[476] +7 * image_in[477] +11 * image_in[478] +41 * image_in[479]
                            +22 * image_in[480] -10 * image_in[481] -32 * image_in[482] -37 * image_in[483] -45 * image_in[484] -45 * image_in[485] -33 * image_in[486] -11 * image_in[487] +2 * image_in[488] +1 * image_in[489] -17 * image_in[490] -11 * image_in[491] +6 * image_in[492] +22 * image_in[493] +28 * image_in[494] +27 * image_in[495] +8 * image_in[496] +22 * image_in[497] +23 * image_in[498] +45 * image_in[499] +19 * image_in[500] -31 * image_in[501] +32 * image_in[502] -2 * image_in[503] +12 * image_in[505] +8 * image_in[506] +62 * image_in[507] +14 * image_in[508] +12 * image_in[509] +7 * image_in[510] -21 * image_in[511]
                            -34 * image_in[512] -34 * image_in[513] -36 * image_in[514] -22 * image_in[515] +3 * image_in[516] -4 * image_in[517] -15 * image_in[518] +5 * image_in[519] +22 * image_in[520] +31 * image_in[521] +23 * image_in[522] +30 * image_in[523] +22 * image_in[524] +17 * image_in[525] +53 * image_in[526] +48 * image_in[527] +48 * image_in[528] +10 * image_in[529] -16 * image_in[530] -7 * image_in[531] +4 * image_in[532] +5 * image_in[533] +4 * image_in[534] +37 * image_in[535] +45 * image_in[536] +36 * image_in[537] +15 * image_in[538] +16 * image_in[539] +13 * image_in[540] +7 * image_in[541] -2 * image_in[542] -25 * image_in[543]
                            -8 * image_in[544] +4 * image_in[546] +24 * image_in[547] +22 * image_in[548] +31 * image_in[549] +42 * image_in[550] +30 * image_in[551] +16 * image_in[552] +32 * image_in[553] +41 * image_in[554] +62 * image_in[555] +15 * image_in[556] -29 * image_in[557] -48 * image_in[558] -17 * image_in[559] +2 * image_in[560] -4 * image_in[561] -3 * image_in[562] +42 * image_in[563] +25 * image_in[564] +34 * image_in[565] +29 * image_in[566] +28 * image_in[567] +29 * image_in[568] +26 * image_in[569] +22 * image_in[570] -7 * image_in[571] -2 * image_in[572] +9 * image_in[573] +20 * image_in[575]
                            +12 * image_in[576] +27 * image_in[577] +30 * image_in[578] +29 * image_in[579] +35 * image_in[580] +37 * image_in[581] +48 * image_in[582] +38 * image_in[583] -5 * image_in[584] +5 * image_in[585] -23 * image_in[586] -2 * image_in[587] -6 * image_in[588] +7 * image_in[589] +3 * image_in[590] +31 * image_in[591] +22 * image_in[592] +14 * image_in[593] +25 * image_in[594] +23 * image_in[595] +27 * image_in[596] +18 * image_in[597] +11 * image_in[598] +13 * image_in[599] +17 * image_in[600] +30 * image_in[601] +19 * image_in[602] +16 * image_in[603] +15 * image_in[604] +25 * image_in[605] +23 * image_in[606] +33 * image_in[607]
                            +24 * image_in[608] +30 * image_in[609] +45 * image_in[610] +18 * image_in[611] -30 * image_in[612] -4 * image_in[613] -15 * image_in[614] -5 * image_in[615] +5 * image_in[616] +6 * image_in[617] +23 * image_in[618] +25 * image_in[619] +28 * image_in[620] -14 * image_in[621] -7 * image_in[622] +15 * image_in[623] -10 * image_in[624] +1 * image_in[625] -1 * image_in[626] +15 * image_in[627] +22 * image_in[628] +17 * image_in[629] +14 * image_in[630] +22 * image_in[631] +14 * image_in[632] +16 * image_in[633] +32 * image_in[634] +9 * image_in[635] +31 * image_in[636] +21 * image_in[637] +21 * image_in[638] -8 * image_in[639]
                            -24 * image_in[640] -7 * image_in[641] -14 * image_in[642] +3 * image_in[643] +6 * image_in[644] -4 * image_in[645] +21 * image_in[646] +59 * image_in[647] +47 * image_in[648] +12 * image_in[649] -1 * image_in[650] +13 * image_in[651] +21 * image_in[652] +19 * image_in[653] +13 * image_in[654] +4 * image_in[655] +3 * image_in[656] +7 * image_in[657] +7 * image_in[658] +19 * image_in[659] +20 * image_in[660] +6 * image_in[661] +10 * image_in[662] +32 * image_in[663] +34 * image_in[664] -10 * image_in[665] +6 * image_in[666] +2 * image_in[667] +4 * image_in[668] -3 * image_in[669] -19 * image_in[670] -1 * image_in[671]
                            -3 * image_in[672] +3 * image_in[673] +15 * image_in[674] +36 * image_in[675] +27 * image_in[676] -13 * image_in[677] +12 * image_in[678] +33 * image_in[679] +17 * image_in[680] +30 * image_in[681] +13 * image_in[682] +36 * image_in[683] +28 * image_in[684] +33 * image_in[685] +41 * image_in[686] +35 * image_in[687] +36 * image_in[688] +18 * image_in[689] +20 * image_in[690] +23 * image_in[691] -10 * image_in[692] +10 * image_in[693] -6 * image_in[694] +1 * image_in[695] +15 * image_in[696] +14 * image_in[697] +5 * image_in[698] +6 * image_in[699] -6 * image_in[701] -4 * image_in[702] +9 * image_in[703]
                            -2 * image_in[704] -1 * image_in[705] +28 * image_in[706] +26 * image_in[707] +44 * image_in[708] +42 * image_in[709] +52 * image_in[710] +41 * image_in[711] +63 * image_in[712] +37 * image_in[713] +36 * image_in[714] +36 * image_in[715] +41 * image_in[716] +30 * image_in[717] +12 * image_in[718] +20 * image_in[719] -1 * image_in[720] +2 * image_in[721] +38 * image_in[722] +15 * image_in[723] +19 * image_in[724] +2 * image_in[725] +2 * image_in[726] -4 * image_in[727] +5 * image_in[728] +5 * image_in[730] +2 * image_in[731] -13 * image_in[732] -22 * image_in[733] -4 * image_in[734] -10 * image_in[735]
                            -19 * image_in[736] +7 * image_in[737] -10 * image_in[738] +4 * image_in[740] +1 * image_in[741] -24 * image_in[742] +2 * image_in[743] -6 * image_in[744] -17 * image_in[745] -12 * image_in[746] -23 * image_in[747] -8 * image_in[748] -3 * image_in[749] +5 * image_in[750] +7 * image_in[751] +4 * image_in[752] -5 * image_in[753] -6 * image_in[755] -5 * image_in[756] +3 * image_in[757] +1 * image_in[758] +5 * image_in[759] +1 * image_in[760] -8 * image_in[761] -17 * image_in[762] -30 * image_in[763] -30 * image_in[764] -30 * image_in[765] -29 * image_in[766] +13 * image_in[767]
                            +9 * image_in[768] -39 * image_in[769] -23 * image_in[770] -23 * image_in[771] -41 * image_in[772] -53 * image_in[773] -32 * image_in[774] -19 * image_in[775] -40 * image_in[776] -21 * image_in[777] -6 * image_in[778] -2 * image_in[779] -4 * image_in[780] -5 * image_in[781] -3 * image_in[782] +2 * image_in[783];
                        if (layer1_out[15] < 0) layer1_out[15] = 0;
                        counter <= counter + 1;
                    end else begin
                        state <= LAYER2;
                        counter <= 0;
                    end
                end

                LAYER2: begin
                    // 计算第二层（10个神经元）
                    if (counter == 0) begin
                        layer2_out[0] = -99 - ((19 * layer1_out[0]) >>> 7) + ((11 * layer1_out[1]) >>> 7) - ((44 * layer1_out[2]) >>> 7) + ((33 * layer1_out[3]) >>> 7) - ((73 * layer1_out[4]) >>> 7) + ((36 * layer1_out[5]) >>> 7) + ((37 * layer1_out[6]) >>> 7) + ((53 * layer1_out[7]) >>> 7) + ((16 * layer1_out[8]) >>> 7) + ((58 * layer1_out[9]) >>> 7) - ((13 * layer1_out[10]) >>> 7) - ((64 * layer1_out[11]) >>> 7) - ((105 * layer1_out[12]) >>> 7) + ((8 * layer1_out[13]) >>> 7) - ((43 * layer1_out[14]) >>> 7) - ((70 * layer1_out[15]) >>> 7);
                        layer2_out[1] = 66 + ((31 * layer1_out[0]) >>> 7) - ((9 * layer1_out[1]) >>> 7) - ((65 * layer1_out[2]) >>> 7) - ((118 * layer1_out[3]) >>> 7) + ((62 * layer1_out[4]) >>> 7) - ((21 * layer1_out[5]) >>> 7) - ((94 * layer1_out[6]) >>> 7) - ((36 * layer1_out[7]) >>> 7) - ((121 * layer1_out[8]) >>> 7) + ((78 * layer1_out[9]) >>> 7) + ((67 * layer1_out[10]) >>> 7) - ((54 * layer1_out[11]) >>> 7) + ((48 * layer1_out[12]) >>> 7) + ((23 * layer1_out[13]) >>> 7) - ((13 * layer1_out[14]) >>> 7) - ((14 * layer1_out[15]) >>> 7);
                        layer2_out[2] = -5 + ((23 * layer1_out[0]) >>> 7) + ((41 * layer1_out[1]) >>> 7) - ((69 * layer1_out[2]) >>> 7) + ((35 * layer1_out[3]) >>> 7) + ((20 * layer1_out[4]) >>> 7) + ((31 * layer1_out[5]) >>> 7) - ((39 * layer1_out[6]) >>> 7) + ((3 * layer1_out[7]) >>> 7) + ((44 * layer1_out[8]) >>> 7) - ((68 * layer1_out[9]) >>> 7) - ((102 * layer1_out[10]) >>> 7) + ((45 * layer1_out[11]) >>> 7) + ((10 * layer1_out[12]) >>> 7) + ((4 * layer1_out[13]) >>> 7) - ((27 * layer1_out[14]) >>> 7) + ((1 * layer1_out[15]) >>> 7);
                        layer2_out[3] = 27 - ((31 * layer1_out[0]) >>> 7) + ((66 * layer1_out[1]) >>> 7) - ((9 * layer1_out[2]) >>> 7) - ((34 * layer1_out[3]) >>> 7) + ((35 * layer1_out[4]) >>> 7) - ((2 * layer1_out[5]) >>> 7) + ((50 * layer1_out[6]) >>> 7) - ((87 * layer1_out[7]) >>> 7) - ((36 * layer1_out[8]) >>> 7) + ((20 * layer1_out[9]) >>> 7) - ((29 * layer1_out[10]) >>> 7) - ((43 * layer1_out[11]) >>> 7) - ((27 * layer1_out[12]) >>> 7) - ((36 * layer1_out[13]) >>> 7) - ((84 * layer1_out[14]) >>> 7) + ((52 * layer1_out[15]) >>> 7);
                        layer2_out[4] = 10 + ((9 * layer1_out[0]) >>> 7) - ((127 * layer1_out[1]) >>> 7) + ((43 * layer1_out[2]) >>> 7) - ((36 * layer1_out[3]) >>> 7) + ((36 * layer1_out[4]) >>> 7) - ((93 * layer1_out[5]) >>> 7) + ((34 * layer1_out[6]) >>> 7) + ((5 * layer1_out[7]) >>> 7) + ((19 * layer1_out[8]) >>> 7) - ((78 * layer1_out[9]) >>> 7) - ((47 * layer1_out[10]) >>> 7) - ((34 * layer1_out[11]) >>> 7) - ((90 * layer1_out[12]) >>> 7) + ((68 * layer1_out[13]) >>> 7) - ((1 * layer1_out[14]) >>> 7) - ((62 * layer1_out[15]) >>> 7);
                        layer2_out[5] = 127 + ((53 * layer1_out[0]) >>> 7) - ((37 * layer1_out[1]) >>> 7) - ((22 * layer1_out[2]) >>> 7) - ((52 * layer1_out[3]) >>> 7) - ((31 * layer1_out[4]) >>> 7) - ((27 * layer1_out[5]) >>> 7) + ((60 * layer1_out[6]) >>> 7) + ((53 * layer1_out[7]) >>> 7) - ((22 * layer1_out[8]) >>> 7) + ((36 * layer1_out[9]) >>> 7) - ((22 * layer1_out[10]) >>> 7) - ((75 * layer1_out[11]) >>> 7) + ((16 * layer1_out[12]) >>> 7) - ((44 * layer1_out[13]) >>> 7) - ((13 * layer1_out[14]) >>> 7) + ((48 * layer1_out[15]) >>> 7);
                        layer2_out[6] = -16 - ((55 * layer1_out[0]) >>> 7) - ((73 * layer1_out[1]) >>> 7) - ((35 * layer1_out[2]) >>> 7) - ((71 * layer1_out[3]) >>> 7) + ((18 * layer1_out[4]) >>> 7) + ((16 * layer1_out[5]) >>> 7) - ((20 * layer1_out[6]) >>> 7) + ((44 * layer1_out[7]) >>> 7) + ((59 * layer1_out[8]) >>> 7) + ((14 * layer1_out[9]) >>> 7) - ((24 * layer1_out[10]) >>> 7) + ((68 * layer1_out[11]) >>> 7) - ((69 * layer1_out[12]) >>> 7) + ((6 * layer1_out[13]) >>> 7) + ((71 * layer1_out[14]) >>> 7) - ((3 * layer1_out[15]) >>> 7);
                        layer2_out[7] = 12 - ((59 * layer1_out[0]) >>> 7) + ((5 * layer1_out[1]) >>> 7) + ((40 * layer1_out[2]) >>> 7) + ((34 * layer1_out[3]) >>> 7) - ((30 * layer1_out[4]) >>> 7) - ((69 * layer1_out[5]) >>> 7) + ((24 * layer1_out[6]) >>> 7) - ((16 * layer1_out[7]) >>> 7) - ((53 * layer1_out[8]) >>> 7) + ((59 * layer1_out[9]) >>> 7) + ((3 * layer1_out[10]) >>> 7) + ((71 * layer1_out[11]) >>> 7) + ((66 * layer1_out[12]) >>> 7) + ((37 * layer1_out[13]) >>> 7) - ((95 * layer1_out[14]) >>> 7) - ((61 * layer1_out[15]) >>> 7);
                        layer2_out[8] = -85 + ((43 * layer1_out[0]) >>> 7) - ((16 * layer1_out[1]) >>> 7) + ((25 * layer1_out[2]) >>> 7) + ((8 * layer1_out[3]) >>> 7) - ((46 * layer1_out[4]) >>> 7) + ((10 * layer1_out[5]) >>> 7) - ((3 * layer1_out[6]) >>> 7) - ((58 * layer1_out[7]) >>> 7) - ((74 * layer1_out[8]) >>> 7) - ((89 * layer1_out[9]) >>> 7) + ((3 * layer1_out[10]) >>> 7) - ((29 * layer1_out[11]) >>> 7) - ((55 * layer1_out[12]) >>> 7) + ((17 * layer1_out[13]) >>> 7) + ((40 * layer1_out[14]) >>> 7) + ((36 * layer1_out[15]) >>> 7);
                        layer2_out[9] = -20 - ((29 * layer1_out[0]) >>> 7) - ((76 * layer1_out[1]) >>> 7) + ((60 * layer1_out[2]) >>> 7) + ((71 * layer1_out[3]) >>> 7) + ((24 * layer1_out[4]) >>> 7) - ((41 * layer1_out[5]) >>> 7) + ((10 * layer1_out[6]) >>> 7) - ((41 * layer1_out[7]) >>> 7) + ((5 * layer1_out[8]) >>> 7) - ((51 * layer1_out[9]) >>> 7) + ((27 * layer1_out[10]) >>> 7) - ((96 * layer1_out[11]) >>> 7) - ((1 * layer1_out[12]) >>> 7) - ((74 * layer1_out[13]) >>> 7) - ((7 * layer1_out[14]) >>> 7) - ((45 * layer1_out[15]) >>> 7);
                        counter <= counter + 1;
                    end else begin
                        state <= DONE;
                    end
                end

                DONE: begin
                    // 找到最大值的索引
                    if (layer2_out[0] >= layer2_out[1] && layer2_out[0] >= layer2_out[2] &&
                        layer2_out[0] >= layer2_out[3] && layer2_out[0] >= layer2_out[4] &&
                        layer2_out[0] >= layer2_out[5] && layer2_out[0] >= layer2_out[6] &&
                        layer2_out[0] >= layer2_out[7] && layer2_out[0] >= layer2_out[8] &&
                        layer2_out[0] >= layer2_out[9])
                        digit_out <= 0;
                    else if (layer2_out[1] >= layer2_out[2] && layer2_out[1] >= layer2_out[3] &&
                             layer2_out[1] >= layer2_out[4] && layer2_out[1] >= layer2_out[5] &&
                             layer2_out[1] >= layer2_out[6] && layer2_out[1] >= layer2_out[7] &&
                             layer2_out[1] >= layer2_out[8] && layer2_out[1] >= layer2_out[9])
                        digit_out <= 1;
                    else if (layer2_out[2] >= layer2_out[3] && layer2_out[2] >= layer2_out[4] &&
                             layer2_out[2] >= layer2_out[5] && layer2_out[2] >= layer2_out[6] &&
                             layer2_out[2] >= layer2_out[7] && layer2_out[2] >= layer2_out[8] &&
                             layer2_out[2] >= layer2_out[9])
                        digit_out <= 2;
                    else if (layer2_out[3] >= layer2_out[4] && layer2_out[3] >= layer2_out[5] &&
                             layer2_out[3] >= layer2_out[6] && layer2_out[3] >= layer2_out[7] &&
                             layer2_out[3] >= layer2_out[8] && layer2_out[3] >= layer2_out[9])
                        digit_out <= 3;
                    else if (layer2_out[4] >= layer2_out[5] && layer2_out[4] >= layer2_out[6] &&
                             layer2_out[4] >= layer2_out[7] && layer2_out[4] >= layer2_out[8] &&
                             layer2_out[4] >= layer2_out[9])
                        digit_out <= 4;
                    else if (layer2_out[5] >= layer2_out[6] && layer2_out[5] >= layer2_out[7] &&
                             layer2_out[5] >= layer2_out[8] && layer2_out[5] >= layer2_out[9])
                        digit_out <= 5;
                    else if (layer2_out[6] >= layer2_out[7] && layer2_out[6] >= layer2_out[8] &&
                             layer2_out[6] >= layer2_out[9])
                        digit_out <= 6;
                    else if (layer2_out[7] >= layer2_out[8] && layer2_out[7] >= layer2_out[9])
                        digit_out <= 7;
                    else if (layer2_out[8] >= layer2_out[9])
                        digit_out <= 8;
                    else
                        digit_out <= 9;

                    valid <= 1;
                    state <= IDLE;
                end
            endcase
        end
    end

endmodule
